//---Example Use---
// charizard image1 (
//	.pixel(),
//	.color(),
//	.width(),
//	.height()
//);

module charizard (
	input wire [16:0] pixel,
	output wire [8:0] width, height,
	output reg [15:0] color
);

	reg [15:0] image [3248:0] = '{
		16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff,
		16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'h1882, 16'h1882, 16'h1882, 16'h1882, 16'h1882, 16'h1882, 16'h1882, 16'h1882, 16'h1882, 16'h1882, 16'h1882, 16'h1882, 16'h1882, 16'h1882, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff,
		16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'h1882, 16'h1882, 16'h1882, 16'h1882, 16'h1882, 16'h1882, 16'h1882, 16'h1882, 16'h1882, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'h1882, 16'h1882, 16'h1882, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff,
		16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'h1882, 16'h1882, 16'h1882, 16'h1882, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'h1882, 16'h1882, 16'h1882, 16'h1882, 16'h1882, 16'h1882, 16'h1882, 16'h1882, 16'h1882, 16'h1882, 16'h1882, 16'h1882, 16'h1882, 16'h1882, 16'h1882, 16'h1882, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff,
		16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'h1882, 16'h1882, 16'h1882, 16'hf5a, 16'hf5a, 16'hf5a, 16'h1882, 16'h1882, 16'hf5a, 16'hf5a, 16'hf5a, 16'hd286, 16'hd286, 16'h1882, 16'h1882, 16'h1882, 16'h1882, 16'h1882, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hf5a, 16'hf5a, 16'hf5a, 16'h1882, 16'h1882, 16'h1882, 16'h1882, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff,
		16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'h1882, 16'h1882, 16'hffff, 16'hd286, 16'hf5a, 16'hf5a, 16'hf5a, 16'h1882, 16'hd286, 16'hffff, 16'h1882, 16'h1882, 16'h1882, 16'h1882, 16'h1882, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'hf5a, 16'hf5a, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hf5a, 16'hf5a, 16'hf5a, 16'h1882, 16'h1882, 16'h1882, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff,
		16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'h1882, 16'hffff, 16'hffff, 16'hf5a, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'h1882, 16'hf5a, 16'hffff, 16'h1882, 16'h1882, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'hf5a, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hf5a, 16'h1882, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff,
		16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'h1882, 16'h1882, 16'h1882, 16'h1882, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'h1882, 16'hf5a, 16'hffff, 16'h1882, 16'h1882, 16'h1882, 16'h1882, 16'h1882, 16'h1882, 16'h1882, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'hffff, 16'hffff, 16'hffff, 16'h1882, 16'hd286, 16'h1882, 16'h1882, 16'h1882, 16'h1882, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff,
		16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'h1882, 16'h1882, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'h1882, 16'hf5a, 16'hffff, 16'h1882, 16'h1882, 16'hd286, 16'hf5a, 16'hf5a, 16'hd286, 16'h1882, 16'h1882, 16'h1882, 16'hf5a, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hd286, 16'hd286, 16'hffff, 16'h1882, 16'h1882, 16'hd286, 16'hd286, 16'hf5a, 16'h1882, 16'hd286, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hd286, 16'h1882, 16'hffff, 16'hffff,
		16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'h1882, 16'h1882, 16'h1882, 16'hd286, 16'hd286, 16'h1882, 16'hf5a, 16'hf5a, 16'h1882, 16'h1882, 16'hf5a, 16'hffff, 16'hffff, 16'hffff, 16'h1882, 16'hf5a, 16'h1882, 16'hf5a, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hd286, 16'hd286, 16'hf5a, 16'h1882, 16'h1882, 16'h1882, 16'h1882, 16'h1882, 16'h1882, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hd286, 16'hffff, 16'hffff, 16'hd286, 16'hffff,
		16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'h1882, 16'h1882, 16'h1882, 16'h1882, 16'hd286, 16'hf5a, 16'hf5a, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'h1882, 16'hf5a, 16'hffff, 16'h1882, 16'hf5a, 16'hf5a, 16'hf5a, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'h1882, 16'hf5a, 16'hf5a, 16'hf5a, 16'h1882, 16'hd286, 16'hf5a, 16'hf5a, 16'h1882, 16'h1882, 16'hd286, 16'hffff, 16'hffff, 16'hffff, 16'hd286, 16'h1882, 16'hf5a, 16'h1882, 16'h1882, 16'hffff,
		16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'h1882, 16'h1882, 16'h1882, 16'h1882, 16'h1882, 16'hd286, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'h1882, 16'h1882, 16'hffff, 16'h1882, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'h1882, 16'h1882, 16'hf5a, 16'hf5a, 16'hf5a, 16'hd286, 16'hd286, 16'h1882, 16'hd286, 16'h1882, 16'hffff, 16'hffff, 16'hffff, 16'h1882, 16'hffff, 16'hffff, 16'h1882, 16'h1882, 16'h1882, 16'hffff, 16'h1882, 16'hffff,
		16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'h1882, 16'h1882, 16'h1882, 16'h1882, 16'hd286, 16'hf5a, 16'hf5a, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'h1882, 16'hd286, 16'h1882, 16'hf5a, 16'h1882, 16'hf5a, 16'hf5a, 16'h1882, 16'h1882, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'h1882, 16'h1882, 16'hd286, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'h1882, 16'hffff, 16'h1882, 16'hffff, 16'h1882, 16'hf5a, 16'h1882, 16'hffff,
		16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'h1882, 16'hd286, 16'h1882, 16'hd286, 16'hf5a, 16'hf5a, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'h1882, 16'hf5a, 16'hf5a, 16'hf5a, 16'hd286, 16'h1882, 16'h1882, 16'h1882, 16'h1882, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'h1882, 16'h1882, 16'hd286, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hffff, 16'hffff, 16'h1882, 16'h1882, 16'hffff, 16'h1882, 16'hf5a, 16'h1882, 16'hffff,
		16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'h1882, 16'hd286, 16'hd286, 16'h1882, 16'hd286, 16'hf5a, 16'hf5a, 16'hf5a, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hf5a, 16'hf5a, 16'hf5a, 16'hffff, 16'hf5a, 16'hf5a, 16'hffff, 16'hffff, 16'hffff, 16'hd286, 16'h1882, 16'h1882, 16'h1882, 16'h1882, 16'hd286, 16'hd286, 16'h1882, 16'h1882, 16'h1882, 16'hd286, 16'hd286, 16'hd286, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hffff, 16'h1882, 16'hffff, 16'h1882, 16'hf5a, 16'h1882, 16'hffff,
		16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'h1882, 16'hd286, 16'hd286, 16'h1882, 16'hd286, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hffff, 16'hffff, 16'hf5a, 16'hd286, 16'hd286, 16'hd286, 16'hf5a, 16'hffff, 16'hf5a, 16'hf5a, 16'hffff, 16'hffff, 16'hffff, 16'hf5a, 16'h1882, 16'h1882, 16'h1882, 16'h1882, 16'h1882, 16'h1882, 16'h1882, 16'h1882, 16'h1882, 16'hd286, 16'hd286, 16'hd286, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hd286, 16'hf5a, 16'hffff, 16'h1882, 16'h1882, 16'hffff,
		16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'h1882, 16'h1882, 16'h1882, 16'h1882, 16'h1882, 16'h1882, 16'h1882, 16'h1882, 16'hd286, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hd286, 16'hd286, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hd286, 16'hffff, 16'hffff, 16'h1882, 16'h1882, 16'h1882, 16'hd286, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'h1882, 16'h1882, 16'hd286, 16'hd286, 16'hd286, 16'hf5a, 16'hf5a, 16'hf5a, 16'hd286, 16'hf5a, 16'hf5a, 16'hf5a, 16'h1882, 16'hffff,
		16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'h1882, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hd286, 16'hffff, 16'h1882, 16'hd286, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'h1882, 16'hd286, 16'hd286, 16'hd286, 16'hf5a, 16'hf5a, 16'hf5a, 16'hd286, 16'hd286, 16'hd286, 16'h1882, 16'hffff,
		16'hffff, 16'hffff, 16'hffff, 16'h1882, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'h1882, 16'h1882, 16'h1882, 16'h1882, 16'h1882, 16'h1882, 16'h1882, 16'h1882, 16'hd286, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hd286, 16'h1882, 16'h1882, 16'hd286, 16'hd286, 16'hd286, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hffff, 16'h1882, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'h1882, 16'hd286, 16'hd286, 16'hd286, 16'hf5a, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'h1882, 16'hffff,
		16'hffff, 16'hffff, 16'h1882, 16'hffff, 16'h1882, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'h1882, 16'hd286, 16'hd286, 16'hd286, 16'h1882, 16'hd286, 16'hd286, 16'hd286, 16'hf5a, 16'hd286, 16'h1882, 16'h1882, 16'hd286, 16'h1882, 16'hd286, 16'hd286, 16'hd286, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hd286, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'h1882, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'h1882, 16'hffff,
		16'hffff, 16'hffff, 16'h1882, 16'hf5a, 16'hffff, 16'h1882, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'h1882, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'h1882, 16'hd286, 16'hd286, 16'hd286, 16'h1882, 16'hf5a, 16'h1882, 16'h1882, 16'h1882, 16'hd286, 16'hd286, 16'hd286, 16'hf5a, 16'hf5a, 16'hd286, 16'h1882, 16'hf5a, 16'h1882, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hf5a, 16'h1882, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'h1882, 16'h1882, 16'h1882, 16'hffff,
		16'hffff, 16'hffff, 16'h1882, 16'hf5a, 16'hffff, 16'hffff, 16'h1882, 16'h1882, 16'h1882, 16'h1882, 16'h1882, 16'h1882, 16'hd286, 16'h1882, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'h1882, 16'hd286, 16'h1882, 16'hf5a, 16'hffff, 16'hffff, 16'hffff, 16'h1882, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'h1882, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hf5a, 16'h1882, 16'h1882, 16'hd286, 16'hd286, 16'h1882, 16'h1882, 16'hffff, 16'hffff,
		16'hffff, 16'hffff, 16'hffff, 16'h1882, 16'hf5a, 16'hffff, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'h1882, 16'hd286, 16'hd286, 16'hf5a, 16'hf5a, 16'hd286, 16'hd286, 16'h1882, 16'h1882, 16'h1882, 16'h1882, 16'hd286, 16'h1882, 16'h1882, 16'h1882, 16'h1882, 16'hd286, 16'hd286, 16'hd286, 16'h1882, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hf5a, 16'h1882, 16'h1882, 16'h1882, 16'hd286, 16'h1882, 16'hffff, 16'hffff, 16'hffff,
		16'hffff, 16'hffff, 16'hffff, 16'h1882, 16'hf5a, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'h1882, 16'h1882, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'h1882, 16'h1882, 16'h1882, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hf5a, 16'hf5a, 16'h1882, 16'h1882, 16'h1882, 16'hd286, 16'hffff, 16'hffff, 16'hffff,
		16'hffff, 16'hffff, 16'hffff, 16'h1882, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'h1882, 16'h1882, 16'hf5a, 16'hf5a, 16'h1882, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hd286, 16'h1882, 16'hd286, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hf5a, 16'hf5a, 16'h1882, 16'h1882, 16'h1882, 16'hffff, 16'hffff, 16'hffff, 16'hffff,
		16'hffff, 16'hffff, 16'hffff, 16'h1882, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'h1882, 16'h1882, 16'h1882, 16'hd286, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'h1882, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'h1882, 16'hf5a, 16'hffff, 16'hffff, 16'hd286, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hf5a, 16'hf5a, 16'hf5a, 16'h1882, 16'h1882, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff,
		16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'h1882, 16'hd286, 16'h1882, 16'h1882, 16'h1882, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'h1882, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'h1882, 16'hf5a, 16'hf5a, 16'h1882, 16'h1882, 16'hd286, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hf5a, 16'hf5a, 16'hf5a, 16'h1882, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff,
		16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'h1882, 16'hd286, 16'h1882, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hffff, 16'hf5a, 16'h1882, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hd286, 16'hf5a, 16'hd286, 16'h1882, 16'hf5a, 16'hffff, 16'hffff, 16'hd286, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hf5a, 16'hf5a, 16'hf5a, 16'h1882, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff,
		16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'h1882, 16'hd286, 16'hd286, 16'h1882, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hffff, 16'hffff, 16'hf5a, 16'h1882, 16'hf5a, 16'hf5a, 16'hf5a, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'h1882, 16'hf5a, 16'hf5a, 16'hd286, 16'hf5a, 16'hf5a, 16'hf5a, 16'h1882, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hf5a, 16'hf5a, 16'hf5a, 16'hd286, 16'h1882, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff,
		16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'h1882, 16'hd286, 16'hd286, 16'h1882, 16'hd286, 16'hd286, 16'hd286, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hffff, 16'hffff, 16'hf5a, 16'h1882, 16'hf5a, 16'hf5a, 16'hd286, 16'h1882, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'h1882, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hd286, 16'h1882, 16'hd286, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hd286, 16'h1882, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff,
		16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'h1882, 16'hd286, 16'hd286, 16'h1882, 16'hd286, 16'hd286, 16'hd286, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hffff, 16'hffff, 16'hf5a, 16'h1882, 16'hf5a, 16'hffff, 16'hffff, 16'hd286, 16'h1882, 16'hffff, 16'hffff, 16'hffff, 16'h1882, 16'hd286, 16'hf5a, 16'hffff, 16'hf5a, 16'hf5a, 16'hf5a, 16'h1882, 16'hf5a, 16'hffff, 16'h1882, 16'hffff, 16'hd286, 16'h1882, 16'h1882, 16'hd286, 16'hf5a, 16'hf5a, 16'hd286, 16'hd286, 16'h1882, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff,
		16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'h1882, 16'hd286, 16'hd286, 16'h1882, 16'hd286, 16'hd286, 16'hd286, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hffff, 16'hffff, 16'hffff, 16'h1882, 16'hf5a, 16'hf5a, 16'hffff, 16'hffff, 16'hffff, 16'hd286, 16'h1882, 16'hd286, 16'hf5a, 16'hffff, 16'hffff, 16'hffff, 16'hd286, 16'hf5a, 16'hf5a, 16'h1882, 16'hf5a, 16'hf5a, 16'h1882, 16'h1882, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'h1882, 16'hd286, 16'hd286, 16'h1882, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff,
		16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'h1882, 16'hd286, 16'hd286, 16'hd286, 16'h1882, 16'hd286, 16'hd286, 16'hd286, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hffff, 16'hffff, 16'hffff, 16'hf5a, 16'h1882, 16'hf5a, 16'hf5a, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hf5a, 16'hd286, 16'hd286, 16'hf5a, 16'hd286, 16'h1882, 16'hd286, 16'hf5a, 16'hf5a, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hd286, 16'h1882, 16'h1882, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff,
		16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'h1882, 16'hd286, 16'hd286, 16'hd286, 16'h1882, 16'hd286, 16'hd286, 16'hd286, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'h1882, 16'hf5a, 16'hf5a, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hf5a, 16'hd286, 16'hd286, 16'h1882, 16'hd286, 16'hd286, 16'hf5a, 16'hf5a, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'h1882, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff,
		16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'h1882, 16'hd286, 16'hd286, 16'hd286, 16'h1882, 16'hd286, 16'hd286, 16'hd286, 16'hf5a, 16'hf5a, 16'hf5a, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hf5a, 16'h1882, 16'hf5a, 16'hf5a, 16'hf5a, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hf5a, 16'hf5a, 16'hd286, 16'hd286, 16'h1882, 16'hd286, 16'hf5a, 16'hf5a, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hd286, 16'h1882, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff,
		16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'h1882, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'h1882, 16'h1882, 16'hf5a, 16'hd286, 16'hd286, 16'hf5a, 16'hf5a, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'h1882, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hd286, 16'hd286, 16'h1882, 16'hd286, 16'hf5a, 16'hf5a, 16'hf5a, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'h1882, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff,
		16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'h1882, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'h1882, 16'hf5a, 16'hf5a, 16'hd286, 16'hd286, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hf5a, 16'h1882, 16'hd286, 16'hd286, 16'hf5a, 16'hf5a, 16'hf5a, 16'hd286, 16'hd286, 16'hd286, 16'h1882, 16'hd286, 16'hf5a, 16'hf5a, 16'hf5a, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hd286, 16'h1882, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff,
		16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'h1882, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'h1882, 16'hf5a, 16'hf5a, 16'hf5a, 16'hd286, 16'hd286, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hf5a, 16'h1882, 16'h1882, 16'h1882, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'h1882, 16'hd286, 16'hd286, 16'hd286, 16'hf5a, 16'hf5a, 16'hf5a, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'h1882, 16'h1882, 16'hd286, 16'hffff, 16'h1882, 16'h1882, 16'hffff, 16'hffff,
		16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'h1882, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'h1882, 16'h1882, 16'hf5a, 16'hf5a, 16'hf5a, 16'hd286, 16'hd286, 16'hd286, 16'hffff, 16'hffff, 16'hf5a, 16'hf5a, 16'hd286, 16'h1882, 16'h1882, 16'h1882, 16'h1882, 16'h1882, 16'hd286, 16'hd286, 16'hd286, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'h1882, 16'h1882, 16'hffff, 16'hffff, 16'h1882, 16'hffff, 16'hffff, 16'hd286, 16'hffff,
		16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'h1882, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'h1882, 16'h1882, 16'h1882, 16'hf5a, 16'hf5a, 16'hf5a, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'hf5a, 16'hd286, 16'h1882, 16'h1882, 16'h1882, 16'h1882, 16'h1882, 16'hd286, 16'hd286, 16'hd286, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hffff, 16'hffff, 16'hffff, 16'hf5a, 16'hffff, 16'hffff, 16'hffff, 16'h1882, 16'hf5a, 16'hffff, 16'h1882, 16'hffff,
		16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'h1882, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'h1882, 16'h1882, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hd286, 16'hd286, 16'h1882, 16'h1882, 16'h1882, 16'h1882, 16'h1882, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hffff, 16'hf5a, 16'hf5a, 16'hf5a, 16'hffff, 16'hd286, 16'hf5a, 16'hf5a, 16'h1882, 16'hffff,
		16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'h1882, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'h1882, 16'h1882, 16'hf5a, 16'hf5a, 16'hd286, 16'hd286, 16'h1882, 16'h1882, 16'h1882, 16'h1882, 16'hd286, 16'hd286, 16'h1882, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hd286, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'h1882, 16'hf5a, 16'hd286, 16'hffff,
		16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'h1882, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'h1882, 16'h1882, 16'h1882, 16'h1882, 16'h1882, 16'h1882, 16'h1882, 16'hf5a, 16'hd286, 16'hd286, 16'h1882, 16'h1882, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hd286, 16'hd286, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hd286, 16'h1882, 16'hffff, 16'hffff,
		16'hffff, 16'hf5a, 16'hf5a, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hf5a, 16'hf5a, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'h1882, 16'h1882, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'h1882, 16'h1882, 16'h1882, 16'h1882, 16'hf5a, 16'hd286, 16'hd286, 16'hd286, 16'h1882, 16'h1882, 16'h1882, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'hf5a, 16'hd286, 16'h1882, 16'hd286, 16'hf5a, 16'hf5a, 16'hd286, 16'hffff, 16'hffff, 16'hd286, 16'hffff,
		16'hffff, 16'hf5a, 16'hf5a, 16'hf5a, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hf5a, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'h1882, 16'h1882, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'h1882, 16'hf5a, 16'hf5a, 16'hd286, 16'hd286, 16'hd286, 16'h1882, 16'h1882, 16'h1882, 16'h1882, 16'h1882, 16'h1882, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'h1882, 16'h1882, 16'hd286, 16'hd286, 16'hd286, 16'h1882, 16'hf5a, 16'hffff, 16'h1882, 16'hffff,
		16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'h1882, 16'h1882, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'h1882, 16'hf5a, 16'hf5a, 16'hf5a, 16'hd286, 16'hd286, 16'hd286, 16'h1882, 16'h1882, 16'h1882, 16'h1882, 16'h1882, 16'h1882, 16'h1882, 16'h1882, 16'h1882, 16'h1882, 16'h1882, 16'h1882, 16'hd286, 16'hd286, 16'hd286, 16'h1882, 16'hd286, 16'hf5a, 16'h1882, 16'hffff,
		16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hffff, 16'h1882, 16'h1882, 16'h1882, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'h1882, 16'hd286, 16'hf5a, 16'hf5a, 16'hd286, 16'hd286, 16'hd286, 16'h1882, 16'h1882, 16'h1882, 16'h1882, 16'h1882, 16'h1882, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'h1882, 16'hd286, 16'hd286, 16'h1882, 16'h1882, 16'hd286, 16'hd286, 16'hffff,
		16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hf5a, 16'hf5a, 16'hf5a, 16'hffff, 16'hffff, 16'hffff, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hffff, 16'hffff, 16'h1882, 16'h1882, 16'h1882, 16'h1882, 16'hd286, 16'hf5a, 16'hf5a, 16'hf5a, 16'hd286, 16'hd286, 16'hd286, 16'h1882, 16'h1882, 16'h1882, 16'h1882, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'h1882, 16'h1882, 16'hffff, 16'hffff, 16'h1882, 16'hffff, 16'hffff,
		16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'hf5a, 16'hf5a, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'h1882, 16'h1882, 16'h1882, 16'h1882, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'h1882, 16'hf5a, 16'hffff, 16'hffff, 16'hd286, 16'hffff,
		16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'hf5a, 16'hf5a, 16'hd286, 16'hd286, 16'hd286, 16'h1882, 16'h1882, 16'h1882, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hd286, 16'hd286, 16'hf5a, 16'hffff, 16'h1882, 16'hffff,
		16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'h1882, 16'h1882, 16'h1882, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'h1882, 16'hd286, 16'hf5a, 16'hd286, 16'hffff,
		16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'hd286, 16'h1882, 16'h1882, 16'h1882, 16'h1882, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'h1882, 16'hd286, 16'hffff, 16'hffff,
		16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff,
		16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff,
		16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff,
		16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hf5a, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff,
		16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff
};

//	assign width  = 57;
//	assign height = 57;

	assign width  = 56;	//for 0 indexed width
	assign height = 56;	//for 0 indexed Height

	assign color  = image[pixel];

endmodule
