//---Example Use---
// grasstile image1 (
//	.pixel(),
//	.color(),
//	.width(),
//	.height()
//);

module GrassTile (
	input wire [16:0] pixel,
	output wire [8:0] width, height,
	output reg [15:0] color
);

	reg [15:0] image [255:0] = '{
		16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h8673, 16'h96b5, 16'h96b5, 16'h8673, 16'h8673, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5,
		16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h8673, 16'h8673, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h8673, 16'h96b5,
		16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h8673, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5,
		16'h96b5, 16'haef5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'haef5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'haef5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5,
		16'h96b5, 16'haef5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'haef5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5,
		16'h96b5, 16'haef5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h8673, 16'h8673, 16'h96b5, 16'h96b5,
		16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h8673, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h8673, 16'h96b5, 16'h96b5,
		16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h8673, 16'h8673, 16'h96b5,
		16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'haef5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h8673, 16'h96b5,
		16'h8673, 16'h8673, 16'h96b5, 16'h96b5, 16'haef5, 16'h96b5, 16'h8673, 16'h8673, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5,
		16'h96b5, 16'h8673, 16'h8673, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h8673, 16'h8673, 16'h96b5, 16'h96b5, 16'h8673, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5,
		16'h96b5, 16'h96b5, 16'h8673, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h8673, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'haef5, 16'haef5, 16'h96b5,
		16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'haef5, 16'haef5, 16'h96b5,
		16'h96b5, 16'h96b5, 16'h96b5, 16'haef5, 16'haef5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5,
		16'h96b5, 16'h96b5, 16'h96b5, 16'haef5, 16'haef5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h8673, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5,
		16'h96b5, 16'h8673, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'haef5
};

	//assign width  = 16;
	//assign height = 16;

	assign width  = 15;	//for 0 indexed width
	assign height = 15;	//for 0 indexed Height

	assign color  = image[254 - pixel];

endmodule
