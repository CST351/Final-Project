//---Example Use---
// Battle_Scene image1 (
//	.pixel(),
//	.color(),
//	.width(),
//	.height()
//);

module Battle_Scene (
	input wire [16:0] pixel,
	output wire [8:0] width, height,
	output reg [15:0] color
);

	reg [15:0] image [76799:0] = '{
		16'h7b4a, 16'h7b4b, 16'h7b4b, 16'h7b4b, 16'h6ae9, 16'h5a68, 16'h5a88, 16'h6ac9, 16'h73a, 16'h7b4b, 16'h7b4b, 16'h732b, 16'h7b2a, 16'h7b6b, 16'h836b, 16'h8bab, 16'h8bab, 16'h8bab, 16'h8bcc, 16'h93ec, 16'h93ec, 16'h93ed, 16'h94d, 16'h94c, 16'h9cd, 16'h9c2d, 16'h9c2d, 16'h9c2d, 16'ha44e, 16'h9c2e, 16'ha46f, 16'ha48f, 16'ha4b0, 16'ha4b0, 16'hacd0, 16'hacd0, 16'hacd0, 16'h8bec, 16'h3143, 16'h20c1, 16'h18c1, 16'h840, 16'h840, 16'h861, 16'h020, 16'h020, 16'h040, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h040, 16'h040, 16'h040, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h1081, 16'h2923, 16'h2123, 16'h1081, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h18a2, 16'h49e6, 16'h732a, 16'h6267, 16'h5a67, 16'h5a67, 16'h6266, 16'h6267, 16'h6267, 16'h6267, 16'h6267, 16'h6267, 16'h6aa8, 16'h834a, 16'hacaf, 16'h6287, 16'h3143, 16'h020, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h040, 16'h840, 16'h5247, 16'hacb0, 16'hacb0, 16'hacb1, 16'h9c2f, 16'h49a6, 16'h72eb, 16'hac90, 16'hacb0, 16'ha44f, 16'h7b2b, 16'h5a68, 16'h49e7, 16'h6aa9, 16'h93ee, 16'ha46f, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha46f, 16'h93ed, 16'h8bac, 16'h9c2e, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c2e, 16'h9c2e, 16'h9c2f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4e, 16'h9c4f, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9ce, 16'h9ce, 16'h9ce, 16'h9cd, 16'h94d, 16'h94e, 16'h94d, 16'h94d, 16'h94e, 16'h93ee, 16'h94e, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cc, 16'h93cc, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cc, 16'h8bcc, 16'h8bcd, 16'h8bad, 16'h8bcd, 16'h8bad, 16'h8bad, 16'h8bad, 16'h8bac, 16'h8bac, 16'h8b8c, 16'h8bac, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h6ac9, 16'h2924, 16'h20e1, 16'h20c2, 16'h18c1, 16'h18c1, 16'h1061, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h7b4a, 16'h7b2a, 16'h7b2a, 16'h7b2a, 16'h732a, 16'h6aea, 16'h6ae9, 16'h73a, 16'h7b2b, 16'h836b, 16'h7b4b, 16'h732b, 16'h732a, 16'h7b6b, 16'h838c, 16'h8bab, 16'h8bab, 16'h8bab, 16'h8bec, 16'h94d, 16'h94d, 16'h9c2d, 16'h9c2d, 16'h9c2d, 16'h9c2e, 16'h9c4e, 16'ha46d, 16'ha46e, 16'ha46e, 16'h9c4e, 16'ha46f, 16'ha48f, 16'ha490, 16'ha4af, 16'ha4af, 16'hacb0, 16'ha4b0, 16'h8bcc, 16'h3163, 16'h20c1, 16'h18a1, 16'h840, 16'h040, 16'h861, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h040, 16'h040, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h840, 16'h1081, 16'h18a2, 16'h1061, 16'h00, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h00, 16'h1061, 16'h3944, 16'h7b2a, 16'h6267, 16'h5a67, 16'h6267, 16'h5a66, 16'h5a67, 16'h6267, 16'h6267, 16'h6267, 16'h6287, 16'h6aa7, 16'h834a, 16'hacaf, 16'h6288, 16'h3144, 16'h820, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h840, 16'h5a47, 16'hacb0, 16'hb4b1, 16'hacb1, 16'h8bad, 16'h4185, 16'h93cd, 16'hac90, 16'h93ed, 16'h6aea, 16'h49e6, 16'h5a48, 16'h836c, 16'h9c4f, 16'ha46f, 16'ha48f, 16'ha490, 16'ha48f, 16'ha490, 16'ha470, 16'h93ed, 16'h8bac, 16'h9c2e, 16'ha46f, 16'ha46f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9ce, 16'h9ce, 16'h9ce, 16'h9ce, 16'h9ce, 16'h9ce, 16'h94e, 16'h94e, 16'h94e, 16'h94d, 16'h94d, 16'h94d, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93cd, 16'h93ed, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h8bcd, 16'h8bcd, 16'h93ad, 16'h8bcd, 16'h8bcc, 16'h8bcc, 16'h8bad, 16'h8bac, 16'h8bac, 16'h8bac, 16'h8bac, 16'h8b8c, 16'h6ac9, 16'h3123, 16'h20e1, 16'h20c1, 16'h20c1, 16'h20c1, 16'h1061, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h7b4a, 16'h6ae9, 16'h6ae9, 16'h732a, 16'h73a, 16'h73a, 16'h732a, 16'h73a, 16'h6aea, 16'h7b6b, 16'h7b6b, 16'h7b4b, 16'h7b4b, 16'h836b, 16'h838c, 16'h8bac, 16'h8bcb, 16'h8bcb, 16'h93ec, 16'h94c, 16'h94d, 16'h9cd, 16'h9c2c, 16'h9c2c, 16'h9c2d, 16'h9c4e, 16'ha46e, 16'ha46e, 16'ha46f, 16'h9c6f, 16'ha46e, 16'ha48f, 16'ha48f, 16'ha48f, 16'ha4af, 16'ha4b0, 16'ha48f, 16'h8bcc, 16'h2943, 16'h18c1, 16'h18a1, 16'h840, 16'h040, 16'h861, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h040, 16'h040, 16'h040, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h00, 16'h00, 16'h020, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h1081, 16'h3964, 16'h7ba, 16'h6267, 16'h6267, 16'h6267, 16'h5a67, 16'h6267, 16'h6267, 16'h6267, 16'h6267, 16'h6287, 16'h6aa8, 16'h834a, 16'hacaf, 16'h62a7, 16'h3144, 16'h820, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h840, 16'h5a47, 16'hacb0, 16'hb4b1, 16'hacb1, 16'h73a, 16'h49e6, 16'h93ed, 16'h7b2b, 16'h527, 16'h6268, 16'h7b2b, 16'h93cd, 16'h9c2e, 16'ha44f, 16'ha46f, 16'ha46f, 16'ha490, 16'ha490, 16'ha46f, 16'h94e, 16'h8bac, 16'h9c2e, 16'ha46f, 16'ha46f, 16'ha46f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9ce, 16'h9ce, 16'h94e, 16'h94e, 16'h94d, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h93ee, 16'h93ed, 16'h93ee, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h8bcd, 16'h8bcd, 16'h93cc, 16'h93cd, 16'h93cc, 16'h8bcc, 16'h8bac, 16'h8bcc, 16'h8bad, 16'h8bad, 16'h8bac, 16'h8b8c, 16'h6aca, 16'h3143, 16'h20e1, 16'h20c1, 16'h20c1, 16'h18c1, 16'h1060, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h7b4a, 16'h6ae9, 16'h732a, 16'h7b4b, 16'h73a, 16'h73a, 16'h7b2a, 16'h732a, 16'h73a, 16'h836b, 16'h836b, 16'h836b, 16'h836b, 16'h836b, 16'h838c, 16'h8bac, 16'h8bcb, 16'h93cb, 16'h93ec, 16'h93eb, 16'h93ec, 16'h94d, 16'h9cc, 16'h9cc, 16'h9c2c, 16'h9c4d, 16'ha46d, 16'ha46d, 16'ha46e, 16'ha46e, 16'ha46f, 16'ha46f, 16'ha48f, 16'ha48f, 16'ha48f, 16'ha490, 16'ha48f, 16'h8bcd, 16'h2923, 16'h18a2, 16'h10a1, 16'h840, 16'h041, 16'h861, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h040, 16'h040, 16'h040, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h840, 16'h020, 16'h020, 16'h020, 16'h020, 16'h861, 16'h1081, 16'h3984, 16'h73a, 16'h6267, 16'h6267, 16'h6267, 16'h5a67, 16'h5a67, 16'h5a67, 16'h6267, 16'h6267, 16'h6267, 16'h6aa8, 16'h834a, 16'hb4cf, 16'h6aa7, 16'h3143, 16'h820, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h840, 16'h5a67, 16'hacb1, 16'hb4d1, 16'hacb0, 16'h6289, 16'h49c6, 16'h5a48, 16'h5a28, 16'h7b2b, 16'ha44f, 16'ha470, 16'h9c2e, 16'h9c2e, 16'h9c4f, 16'ha44f, 16'ha46f, 16'ha46f, 16'ha46f, 16'h94e, 16'h8bad, 16'h9c2e, 16'ha490, 16'ha490, 16'ha470, 16'ha46f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2f, 16'h9c2e, 16'h9cf, 16'h9c2e, 16'h9c2e, 16'h9ce, 16'h9c2e, 16'h9c2e, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h93ee, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h8bcd, 16'h8bcd, 16'h8bcd, 16'h8bad, 16'h8bad, 16'h8bad, 16'h8bac, 16'h8b8c, 16'h6ae9, 16'h3143, 16'h20e1, 16'h20c2, 16'h20c1, 16'h18c1, 16'h1060, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h7b4a, 16'h62a9, 16'h732a, 16'h7b2a, 16'h7b4b, 16'h7b4b, 16'h7b4b, 16'h7b4b, 16'h7b4b, 16'h836b, 16'h7b6b, 16'h838b, 16'h838b, 16'h836b, 16'h836b, 16'h8bcb, 16'h8bcb, 16'h93cc, 16'h93ec, 16'h93ec, 16'h93ec, 16'h94c, 16'h9c2c, 16'h9c2c, 16'h9c2c, 16'h9c2c, 16'h9c2c, 16'h9c2d, 16'h9c4e, 16'ha44f, 16'ha46f, 16'ha46f, 16'ha48f, 16'ha48f, 16'ha48f, 16'ha48f, 16'h9c6f, 16'h83cd, 16'h2923, 16'h18a1, 16'h10a1, 16'h040, 16'h021, 16'h861, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h040, 16'h040, 16'h040, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h840, 16'h861, 16'h861, 16'h040, 16'h840, 16'h1081, 16'h860, 16'h2924, 16'h72e9, 16'h6267, 16'h5a67, 16'h6267, 16'h6267, 16'h6267, 16'h6267, 16'h6267, 16'h6266, 16'h6267, 16'h6aa8, 16'h834a, 16'hb4f0, 16'h6aa8, 16'h3163, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h040, 16'h840, 16'h5a68, 16'hacd1, 16'hb4d1, 16'hac90, 16'h5a68, 16'h3965, 16'h6289, 16'h94e, 16'hacb0, 16'hacb0, 16'hac90, 16'ha44f, 16'h9c2e, 16'h9c2e, 16'h9c4e, 16'h9c2e, 16'h9c2e, 16'h93ed, 16'h8bcd, 16'h9c2e, 16'ha490, 16'ha490, 16'ha490, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha44f, 16'ha44f, 16'ha450, 16'ha46f, 16'ha46f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h9c4f, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9ce, 16'h9ce, 16'h9ce, 16'h9ce, 16'h94e, 16'h94e, 16'h94d, 16'h94e, 16'h94e, 16'h94e, 16'h94d, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93ed, 16'h93cd, 16'h8bcd, 16'h93cd, 16'h8bcd, 16'h8bcd, 16'h8bad, 16'h8bac, 16'h8bac, 16'h72e9, 16'h3143, 16'h20e1, 16'h20c1, 16'h20c1, 16'h18c1, 16'h1080, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h732a, 16'h6aa9, 16'h73a, 16'h732a, 16'h732a, 16'h7b2b, 16'h7b4b, 16'h7b4b, 16'h7b4b, 16'h7b4b, 16'h7b6b, 16'h7b6c, 16'h836b, 16'h7b6b, 16'h836b, 16'h8bcb, 16'h93eb, 16'h93ec, 16'h94c, 16'h94c, 16'h94c, 16'h94d, 16'h9cd, 16'h9c2d, 16'h9c2d, 16'h9cc, 16'h94b, 16'h9cc, 16'ha44e, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'h9c6f, 16'h9c6f, 16'h9c4f, 16'h83cd, 16'h2923, 16'h18a1, 16'h10a1, 16'h040, 16'h020, 16'h061, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h040, 16'h040, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h860, 16'h1082, 16'h10a1, 16'h040, 16'h861, 16'h861, 16'h040, 16'h213, 16'h72e9, 16'h6267, 16'h5a67, 16'h6267, 16'h6267, 16'h6267, 16'h6266, 16'h6267, 16'h6267, 16'h6267, 16'h6aa8, 16'h834a, 16'hb4f0, 16'h6aa8, 16'h3143, 16'h820, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h040, 16'h840, 16'h5a68, 16'hacd0, 16'hb4d1, 16'ha46f, 16'h5a48, 16'h6aca, 16'ha490, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'ha490, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h94d, 16'h93cc, 16'h8bcd, 16'h9c2e, 16'ha48f, 16'ha490, 16'ha490, 16'ha490, 16'ha46f, 16'ha46f, 16'ha44f, 16'ha46f, 16'ha46f, 16'ha470, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c4e, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4e, 16'h9c4f, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9ce, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94d, 16'h94d, 16'h94e, 16'h93ee, 16'h94e, 16'h93ed, 16'h94d, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ec, 16'h93ed, 16'h93ed, 16'h93cd, 16'h8bcd, 16'h8bcd, 16'h8bcd, 16'h8bcc, 16'h8bac, 16'h72e9, 16'h3143, 16'h20e1, 16'h20c2, 16'h20c1, 16'h18c1, 16'h1080, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h7b4a, 16'h73a, 16'h7b4a, 16'h7b4b, 16'h7b4b, 16'h7b4b, 16'h7b4b, 16'h7b4b, 16'h7b2b, 16'h7b4b, 16'h7b4b, 16'h7b6b, 16'h7b6b, 16'h836b, 16'h838c, 16'h8bab, 16'h8bab, 16'h93cb, 16'h93ec, 16'h93ec, 16'h94c, 16'h93ec, 16'h6ac8, 16'h62a7, 16'h739, 16'h7b49, 16'h838a, 16'h8bcb, 16'h94e, 16'h9c2e, 16'h9c4e, 16'h9c6f, 16'h9c6f, 16'h9c6f, 16'h9c6f, 16'h9c4e, 16'h93ed, 16'h83ab, 16'h2923, 16'h18a1, 16'h10a1, 16'h840, 16'h041, 16'h061, 16'h020, 16'h020, 16'h020, 16'h040, 16'h840, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h040, 16'h040, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h860, 16'h1081, 16'h1081, 16'h040, 16'h1061, 16'h840, 16'h040, 16'h2123, 16'h6ac9, 16'h5a67, 16'h5a68, 16'h6267, 16'h6267, 16'h6267, 16'h6267, 16'h6267, 16'h6267, 16'h6287, 16'h6aa8, 16'h834a, 16'hacaf, 16'h6aa8, 16'h3144, 16'h820, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h040, 16'h840, 16'h5a68, 16'hb4d0, 16'hb4d1, 16'hb4d1, 16'h9c2f, 16'hacb1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hb4d1, 16'hacb1, 16'hacb0, 16'ha470, 16'h9c2f, 16'h9c2e, 16'h94d, 16'h93ed, 16'h9c4f, 16'ha48f, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha44f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9ce, 16'h9ce, 16'h9ce, 16'h9ce, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94d, 16'h94d, 16'h94e, 16'h94e, 16'h93ee, 16'h93ee, 16'h94d, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h8bcd, 16'h8bad, 16'h8bac, 16'h8bac, 16'h72e9, 16'h3143, 16'h20e2, 16'h20c2, 16'h20c1, 16'h18c1, 16'h1080, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h7b4a, 16'h7b4b, 16'h7b4b, 16'h7b4b, 16'h7b4b, 16'h7b6b, 16'h7b6b, 16'h836b, 16'h836c, 16'h836b, 16'h836c, 16'h836c, 16'h836b, 16'h836c, 16'h8bac, 16'h8b8b, 16'h8b8b, 16'h8bab, 16'h93cc, 16'h93cc, 16'h93ec, 16'h8bcb, 16'h41c4, 16'h18a1, 16'h18c1, 16'h211, 16'h2922, 16'h3163, 16'h39a4, 16'h4a5, 16'h5266, 16'h62c8, 16'h6b9, 16'h7b6a, 16'h838b, 16'h8bac, 16'h72ea, 16'h7b4b, 16'h293, 16'h18a1, 16'h1081, 16'h840, 16'h040, 16'h041, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h040, 16'h040, 16'h020, 16'h040, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h860, 16'h860, 16'h860, 16'h861, 16'h861, 16'h020, 16'h040, 16'h2923, 16'h72e9, 16'h6267, 16'h6268, 16'h6267, 16'h6267, 16'h6267, 16'h6267, 16'h6267, 16'h6267, 16'h6288, 16'h6aa8, 16'h834a, 16'hacaf, 16'h62a8, 16'h3164, 16'h820, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h840, 16'h5a68, 16'hb4d1, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacb0, 16'hacb1, 16'ha490, 16'ha46f, 16'ha46f, 16'ha490, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha490, 16'ha470, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9ce, 16'h9ce, 16'h9ce, 16'h9ce, 16'h9ce, 16'h9ce, 16'h94e, 16'h94e, 16'h94d, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94d, 16'h94d, 16'h94d, 16'h93ed, 16'h93ee, 16'h93ee, 16'h93ee, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93ad, 16'h93ad, 16'h8bcc, 16'h72ea, 16'h3144, 16'h20e2, 16'h20c2, 16'h20c1, 16'h20c1, 16'h1080, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h7b4a, 16'h7b4b, 16'h7b4b, 16'h7b4b, 16'h7b6b, 16'h836b, 16'h7b6b, 16'h836b, 16'h836b, 16'h838b, 16'h838b, 16'h838c, 16'h838c, 16'h838c, 16'h8bac, 16'h8bac, 16'h8bab, 16'h8bab, 16'h93cc, 16'h93cc, 16'h93ec, 16'h8bcc, 16'h39a4, 16'h1080, 16'h880, 16'h880, 16'h1080, 16'h1080, 16'h1080, 16'h10a0, 16'h10a1, 16'h10c1, 16'h18c1, 16'h20e2, 16'h2922, 16'h3143, 16'h3985, 16'h732b, 16'h212, 16'h10a1, 16'h1081, 16'h040, 16'h040, 16'h041, 16'h040, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h020, 16'h020, 16'h840, 16'h840, 16'h020, 16'h020, 16'h020, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h860, 16'h840, 16'h840, 16'h861, 16'h820, 16'h020, 16'h040, 16'h2924, 16'h6ae9, 16'h6267, 16'h6267, 16'h6267, 16'h6267, 16'h6267, 16'h6267, 16'h6267, 16'h6268, 16'h6a88, 16'h6aa8, 16'h834a, 16'hac8f, 16'h6287, 16'h3164, 16'h820, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h840, 16'h841, 16'h6268, 16'hb4d1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'ha490, 16'ha490, 16'ha48f, 16'ha46f, 16'ha470, 16'ha490, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4e, 16'h9c2f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9ce, 16'h9ce, 16'h9ce, 16'h9ce, 16'h9ce, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94d, 16'h94d, 16'h94d, 16'h93ee, 16'h93ee, 16'h93ed, 16'h93ed, 16'h93ee, 16'h93ee, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h8bcd, 16'h72ea, 16'h3144, 16'h20e2, 16'h20c1, 16'h20c1, 16'h20c1, 16'h1061, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h7b4a, 16'h7b4a, 16'h7b4b, 16'h7b4b, 16'h7b6b, 16'h836b, 16'h7b6b, 16'h836b, 16'h836c, 16'h838b, 16'h838c, 16'h838c, 16'h83ac, 16'h83ac, 16'h8bcc, 16'h8bcc, 16'h8bcc, 16'h8bcc, 16'h93cc, 16'h93cc, 16'h93ec, 16'h8bcc, 16'h41c5, 16'h1081, 16'h080, 16'h080, 16'h880, 16'h080, 16'h880, 16'h880, 16'h880, 16'h880, 16'h880, 16'h880, 16'h861, 16'h861, 16'h213, 16'h6ba, 16'h20e2, 16'h1080, 16'h880, 16'h020, 16'h040, 16'h840, 16'h020, 16'h040, 16'h040, 16'h040, 16'h020, 16'h020, 16'h040, 16'h040, 16'h020, 16'h040, 16'h040, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h840, 16'h020, 16'h840, 16'h840, 16'h020, 16'h020, 16'h840, 16'h2924, 16'h72c9, 16'h5a67, 16'h6267, 16'h6267, 16'h6267, 16'h6267, 16'h6267, 16'h6267, 16'h6267, 16'h6a87, 16'h72a8, 16'h834a, 16'hac8e, 16'h6287, 16'h3164, 16'h020, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h040, 16'h840, 16'h841, 16'h5a68, 16'hb4d1, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb0, 16'hac90, 16'hacb0, 16'hacb0, 16'hacb0, 16'ha490, 16'hac90, 16'hac90, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha44f, 16'ha46f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4e, 16'h9c4e, 16'h9c2f, 16'h9c2e, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9ce, 16'h9c2e, 16'h9c2e, 16'h9ce, 16'h9ce, 16'h9cd, 16'h9ce, 16'h9ce, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94d, 16'h94e, 16'h94e, 16'h93ee, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ee, 16'h93ed, 16'h93ee, 16'h93ed, 16'h93cd, 16'h93cd, 16'h93cd, 16'h8bcc, 16'h73a, 16'h3144, 16'h20e2, 16'h18e1, 16'h20c1, 16'h20c1, 16'h1080, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h7b2b, 16'h7b4a, 16'h7b4b, 16'h7b4b, 16'h834b, 16'h7b4b, 16'h836b, 16'h836b, 16'h838b, 16'h838c, 16'h838c, 16'h838c, 16'h83ac, 16'h83ac, 16'h8bcc, 16'h8bcb, 16'h8bac, 16'h8bcc, 16'h8bac, 16'h8bac, 16'h8bcc, 16'h8bac, 16'h41a5, 16'h1081, 16'h860, 16'h080, 16'h080, 16'h880, 16'h880, 16'h880, 16'h880, 16'h860, 16'h880, 16'h860, 16'h040, 16'h020, 16'h18c3, 16'h6aea, 16'h20e2, 16'h10a0, 16'h880, 16'h040, 16'h040, 16'h840, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h040, 16'h040, 16'h020, 16'h020, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h020, 16'h840, 16'h020, 16'h020, 16'h020, 16'h840, 16'h3124, 16'h72c9, 16'h6267, 16'h6267, 16'h6267, 16'h6267, 16'h6267, 16'h6267, 16'h6267, 16'h6267, 16'h6a88, 16'h6aa8, 16'h834a, 16'ha46e, 16'h6287, 16'h3164, 16'h820, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h040, 16'h841, 16'h6289, 16'hb4f1, 16'hb4f1, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacb0, 16'ha46f, 16'hacb0, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha48f, 16'ha48f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4e, 16'h9c4f, 16'h9c2f, 16'h9c2e, 16'h9c4e, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9ce, 16'h9ce, 16'h9ce, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h93ed, 16'h93ed, 16'h94d, 16'h94d, 16'h93ee, 16'h94d, 16'h93ed, 16'h93ed, 16'h93ce, 16'h93cd, 16'h93cd, 16'h93cd, 16'h739, 16'h3143, 16'h20e2, 16'h20e1, 16'h20c1, 16'h20c1, 16'h1080, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h7b2b, 16'h7b4b, 16'h7b4b, 16'h7b4b, 16'h7b6b, 16'h7b6b, 16'h836c, 16'h836b, 16'h838b, 16'h838c, 16'h838c, 16'h838c, 16'h83ac, 16'h83ac, 16'h8bcc, 16'h8bcc, 16'h8bcc, 16'h8bcc, 16'h8bcc, 16'h8bcc, 16'h93cc, 16'h8bcd, 16'h41a5, 16'h1080, 16'h860, 16'h080, 16'h080, 16'h080, 16'h880, 16'h060, 16'h080, 16'h060, 16'h060, 16'h080, 16'h040, 16'h040, 16'h20e3, 16'h62ca, 16'h20c2, 16'h1081, 16'h860, 16'h020, 16'h040, 16'h040, 16'h040, 16'h040, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h040, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h020, 16'h00, 16'h00, 16'h00, 16'h820, 16'h3164, 16'h72e9, 16'h5a67, 16'h6267, 16'h6267, 16'h6267, 16'h6267, 16'h6267, 16'h6267, 16'h6267, 16'h6287, 16'h6aa8, 16'h834a, 16'ha46e, 16'h6287, 16'h3144, 16'h820, 16'h020, 16'h00, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h040, 16'h040, 16'h861, 16'h6289, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacb0, 16'ha490, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9ce, 16'h9ce, 16'h9ce, 16'h9ce, 16'h9c2e, 16'h9ce, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h93ed, 16'h94e, 16'h94e, 16'h94d, 16'h94e, 16'h94d, 16'h94d, 16'h93ee, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93cd, 16'h73a, 16'h3143, 16'h20e2, 16'h18e1, 16'h20c1, 16'h18c1, 16'h1080, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h7b2a, 16'h7b2a, 16'h7b4b, 16'h7b4b, 16'h7b6b, 16'h7b6b, 16'h836b, 16'h836b, 16'h838b, 16'h838c, 16'h838c, 16'h838c, 16'h83ac, 16'h8bac, 16'h8bcc, 16'h8bcd, 16'h8bcc, 16'h8bec, 16'h93ec, 16'h8bcc, 16'h93ec, 16'h8bec, 16'h41c5, 16'h1080, 16'h860, 16'h860, 16'h880, 16'h080, 16'h080, 16'h060, 16'h060, 16'h060, 16'h060, 16'h060, 16'h040, 16'h040, 16'h20e3, 16'h62c9, 16'h20c2, 16'h1081, 16'h860, 16'h020, 16'h040, 16'h040, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h040, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h00, 16'h00, 16'h00, 16'h820, 16'h3964, 16'h6ae9, 16'h5a67, 16'h5a67, 16'h6267, 16'h6267, 16'h6267, 16'h6267, 16'h6267, 16'h6287, 16'h6287, 16'h6aa8, 16'h8349, 16'ha44d, 16'h6287, 16'h3164, 16'h820, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h040, 16'h040, 16'h841, 16'h6289, 16'hb4f1, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hb4d1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb1, 16'hacb0, 16'hacb0, 16'hac90, 16'ha490, 16'ha490, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha48f, 16'ha48f, 16'ha470, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4e, 16'h9c4e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9ce, 16'h9ce, 16'h9ce, 16'h9c2e, 16'h9c2e, 16'h94e, 16'h94e, 16'h9ce, 16'h9ce, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94d, 16'h94e, 16'h94d, 16'h94d, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93cd, 16'h73a, 16'h3143, 16'h20e1, 16'h18e1, 16'h20c1, 16'h18c1, 16'h1080, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h73a, 16'h732a, 16'h7b4a, 16'h7b4b, 16'h836b, 16'h836b, 16'h836b, 16'h836b, 16'h838b, 16'h838b, 16'h838c, 16'h83ac, 16'h83ab, 16'h83cc, 16'h8bcc, 16'h94d, 16'h94d, 16'h94d, 16'h94d, 16'h94d, 16'h94d, 16'h94d, 16'h41e5, 16'h10a0, 16'h060, 16'h860, 16'h860, 16'h080, 16'h080, 16'h060, 16'h080, 16'h080, 16'h060, 16'h060, 16'h040, 16'h040, 16'h213, 16'h62c9, 16'h18c2, 16'h1081, 16'h860, 16'h020, 16'h040, 16'h040, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h020, 16'h040, 16'h020, 16'h020, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h00, 16'h00, 16'h00, 16'h840, 16'h3964, 16'h72c9, 16'h5a47, 16'h6267, 16'h6267, 16'h5a67, 16'h6267, 16'h6267, 16'h6267, 16'h6267, 16'h6287, 16'h6aa8, 16'h834a, 16'h9c4e, 16'h6267, 16'h3163, 16'h020, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h040, 16'h040, 16'h861, 16'h6289, 16'hb4f1, 16'hb4f2, 16'hb512, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hacb0, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha48f, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha44f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c4e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9ce, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9ce, 16'h94e, 16'h9ce, 16'h9c2e, 16'h94e, 16'h94e, 16'h94e, 16'h9ce, 16'h94e, 16'h94e, 16'h93ed, 16'h94d, 16'h93ee, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93cd, 16'h73a, 16'h3144, 16'h20e2, 16'h20c1, 16'h20c1, 16'h18c1, 16'h1081, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h5246, 16'h5a88, 16'h6ae9, 16'h7b4a, 16'h7b4b, 16'h7b6b, 16'h836b, 16'h836b, 16'h838b, 16'h838b, 16'h838c, 16'h83ac, 16'h83ab, 16'h83cc, 16'h8bcc, 16'h8bec, 16'h8cd, 16'h94d, 16'h942d, 16'h942e, 16'h9c2e, 16'h94d, 16'h41e5, 16'h8a0, 16'h080, 16'h080, 16'h060, 16'h080, 16'h080, 16'h060, 16'h060, 16'h060, 16'h060, 16'h060, 16'h860, 16'h861, 16'h213, 16'h62c9, 16'h18c1, 16'h1081, 16'h860, 16'h020, 16'h020, 16'h040, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h020, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h00, 16'h00, 16'h00, 16'h840, 16'h3964, 16'h72e9, 16'h5a47, 16'h6267, 16'h6267, 16'h6267, 16'h6267, 16'h6267, 16'h6267, 16'h6267, 16'h6a87, 16'h6aa8, 16'h834a, 16'h9c4d, 16'h6267, 16'h3163, 16'h820, 16'h020, 16'h020, 16'h020, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h040, 16'h040, 16'h040, 16'h841, 16'h6289, 16'hb4f2, 16'hb4f2, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd0, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9ce, 16'h9ce, 16'h9c2e, 16'h942e, 16'h942e, 16'h94e, 16'h94e, 16'h9ce, 16'h9ce, 16'h9ce, 16'h94e, 16'h94e, 16'h94d, 16'h93ee, 16'h93ee, 16'h93ed, 16'h93ed, 16'h93ed, 16'h73a, 16'h3144, 16'h20e2, 16'h20c2, 16'h20c1, 16'h18c1, 16'h1080, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h2923, 16'h3144, 16'h5227, 16'h6ac9, 16'h7b4a, 16'h7b6b, 16'h836b, 16'h838b, 16'h838b, 16'h838b, 16'h83ac, 16'h83ac, 16'h83cb, 16'h8bcc, 16'h8bcc, 16'h8bed, 16'h8bed, 16'h94d, 16'h94d, 16'h94e, 16'h942e, 16'h94d, 16'h41e5, 16'h10a0, 16'h060, 16'h060, 16'h060, 16'h060, 16'h860, 16'h060, 16'h060, 16'h060, 16'h060, 16'h860, 16'h20e2, 16'h3184, 16'h3144, 16'h62c9, 16'h18a2, 16'h1081, 16'h861, 16'h020, 16'h040, 16'h040, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h020, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h020, 16'h00, 16'h00, 16'h840, 16'h3965, 16'h72e9, 16'h6267, 16'h6267, 16'h6267, 16'h6267, 16'h6267, 16'h6267, 16'h6267, 16'h6267, 16'h6288, 16'h6aa8, 16'h834a, 16'h9c2d, 16'h6267, 16'h3163, 16'h820, 16'h020, 16'h020, 16'h020, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h040, 16'h040, 16'h840, 16'h860, 16'h6289, 16'hb4f1, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha46f, 16'ha470, 16'ha470, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4e, 16'h9c2f, 16'h9c2f, 16'h9c4e, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h942e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9ce, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94d, 16'h93ed, 16'h93ed, 16'h73a, 16'h3143, 16'h20c2, 16'h20c2, 16'h20c1, 16'h18c1, 16'h1080, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h41a5, 16'h41c6, 16'h5a68, 16'h6ac9, 16'h7b4a, 16'h7b6b, 16'h836b, 16'h838b, 16'h838b, 16'h838b, 16'h83ac, 16'h83ac, 16'h83cb, 16'h8bcc, 16'h8bcc, 16'h8bec, 16'h8cc, 16'h94d, 16'h94d, 16'h942e, 16'h9c2e, 16'h94d, 16'h41e5, 16'h10a0, 16'h060, 16'h060, 16'h060, 16'h060, 16'h060, 16'h060, 16'h060, 16'h060, 16'h060, 16'h060, 16'h18c1, 16'h3184, 16'h3144, 16'h62a9, 16'h18a1, 16'h1081, 16'h860, 16'h020, 16'h020, 16'h040, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h020, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h00, 16'h020, 16'h020, 16'h020, 16'h00, 16'h00, 16'h840, 16'h3964, 16'h72e9, 16'h6267, 16'h6267, 16'h6267, 16'h6267, 16'h6267, 16'h6267, 16'h6268, 16'h6268, 16'h6288, 16'h6aa8, 16'h834a, 16'h9c2d, 16'h6267, 16'h3164, 16'h020, 16'h020, 16'h020, 16'h00, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h040, 16'h040, 16'h840, 16'h861, 16'h6289, 16'hb4f2, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f2, 16'hb4f1, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd0, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha470, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9ce, 16'h9ce, 16'h9ce, 16'h94e, 16'h94d, 16'h94e, 16'h94e, 16'h94d, 16'h93ee, 16'h93ee, 16'h93ed, 16'h73a, 16'h3143, 16'h20e2, 16'h20c1, 16'h20c1, 16'h18c1, 16'h1080, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h6288, 16'h62a9, 16'h72ea, 16'h7b2a, 16'h7b4b, 16'h7b6b, 16'h836b, 16'h836b, 16'h838b, 16'h83ab, 16'h83ac, 16'h83ac, 16'h8bac, 16'h8bcc, 16'h8bec, 16'h8bec, 16'h93ed, 16'h94d, 16'h942e, 16'h942e, 16'h9c2e, 16'h94d, 16'h41e5, 16'h10a1, 16'h860, 16'h860, 16'h860, 16'h060, 16'h860, 16'h060, 16'h060, 16'h060, 16'h060, 16'h060, 16'h040, 16'h860, 16'h213, 16'h5aa8, 16'h18a1, 16'h1081, 16'h860, 16'h020, 16'h040, 16'h040, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h020, 16'h020, 16'h040, 16'h020, 16'h020, 16'h020, 16'h00, 16'h020, 16'h1061, 16'h1082, 16'h1061, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h861, 16'h3164, 16'h72e9, 16'h6267, 16'h6267, 16'h6267, 16'h6267, 16'h6267, 16'h6267, 16'h6267, 16'h6267, 16'h6287, 16'h6aa8, 16'h834a, 16'h9c2d, 16'h6267, 16'h3164, 16'h820, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h040, 16'h840, 16'h860, 16'h6289, 16'hb4f2, 16'hb512, 16'hbd12, 16'hbd12, 16'hbd12, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha470, 16'ha470, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h9c4e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h942e, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h93ed, 16'h732a, 16'h3144, 16'h20e2, 16'h20c1, 16'h20c1, 16'h20c1, 16'h1080, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h73a, 16'h73a, 16'h7b2a, 16'h7b4b, 16'h7b4b, 16'h7b6b, 16'h7b6b, 16'h838b, 16'h838b, 16'h838b, 16'h83ac, 16'h83ac, 16'h8bac, 16'h8bcc, 16'h8bcd, 16'h8bec, 16'h94d, 16'h94d, 16'h942e, 16'h9c2e, 16'h9c2e, 16'h94d, 16'h4a6, 16'h10a1, 16'h060, 16'h060, 16'h860, 16'h060, 16'h860, 16'h860, 16'h060, 16'h060, 16'h060, 16'h060, 16'h040, 16'h040, 16'h213, 16'h5a88, 16'h10a1, 16'h1081, 16'h860, 16'h020, 16'h040, 16'h040, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h020, 16'h020, 16'h040, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h20c3, 16'h3164, 16'h2944, 16'h841, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h1061, 16'h3144, 16'h72ea, 16'h6267, 16'h6267, 16'h6267, 16'h6267, 16'h6267, 16'h6267, 16'h6267, 16'h6267, 16'h6288, 16'h6aa8, 16'h8349, 16'h9cd, 16'h6267, 16'h3163, 16'h820, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h040, 16'h840, 16'h861, 16'h62a9, 16'hb4f2, 16'hb512, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f2, 16'hb4d1, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha48f, 16'ha48f, 16'ha470, 16'ha470, 16'ha46f, 16'ha470, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4e, 16'h9c4e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9ce, 16'h9ce, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h93ed, 16'h7b2b, 16'h3144, 16'h20c3, 16'h20c2, 16'h20c2, 16'h20c1, 16'h1080, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h7b2a, 16'h734a, 16'h7b4b, 16'h7b4b, 16'h7b6b, 16'h7b4b, 16'h7b6b, 16'h838b, 16'h838b, 16'h83ab, 16'h83ab, 16'h83ac, 16'h8bac, 16'h8bcc, 16'h8bcd, 16'h8bed, 16'h94d, 16'h94e, 16'h942e, 16'h9c2e, 16'h9c4f, 16'h94e, 16'h4a6, 16'h10a0, 16'h060, 16'h060, 16'h860, 16'h860, 16'h860, 16'h860, 16'h080, 16'h060, 16'h860, 16'h060, 16'h040, 16'h040, 16'h2923, 16'h5a88, 16'h10a1, 16'h881, 16'h840, 16'h020, 16'h040, 16'h040, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h020, 16'h040, 16'h040, 16'h040, 16'h020, 16'h020, 16'h020, 16'h020, 16'h20e3, 16'h3164, 16'h2943, 16'h840, 16'h020, 16'h020, 16'h020, 16'h020, 16'h821, 16'h18a2, 16'h3144, 16'h72ea, 16'h6247, 16'h6267, 16'h6267, 16'h6267, 16'h6267, 16'h6267, 16'h6267, 16'h6267, 16'h6287, 16'h6aa8, 16'h832a, 16'h9c2d, 16'h5a67, 16'h3164, 16'h820, 16'h020, 16'h020, 16'h020, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h040, 16'h040, 16'h840, 16'h840, 16'h6289, 16'hb4f2, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha44f, 16'ha46f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'ha44f, 16'h9c4f, 16'h9c4e, 16'h9c4e, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9ce, 16'h9ce, 16'h94e, 16'h94e, 16'h94e, 16'h7b2b, 16'h3144, 16'h20c3, 16'h20c2, 16'h20c1, 16'h18c2, 16'h1081, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h732a, 16'h7b2b, 16'h7b4b, 16'h7b4a, 16'h7b6a, 16'h836b, 16'h836b, 16'h838b, 16'h838b, 16'h83ab, 16'h83ac, 16'h83ac, 16'h8bac, 16'h8bcc, 16'h8bcd, 16'h93ed, 16'h94d, 16'h94d, 16'h942e, 16'h9c2e, 16'h9c4e, 16'h942e, 16'h4a6, 16'h1080, 16'h860, 16'h060, 16'h860, 16'h860, 16'h860, 16'h860, 16'h880, 16'h860, 16'h860, 16'h060, 16'h040, 16'h040, 16'h2923, 16'h5268, 16'h1081, 16'h881, 16'h840, 16'h020, 16'h040, 16'h040, 16'h040, 16'h040, 16'h020, 16'h020, 16'h020, 16'h020, 16'h040, 16'h040, 16'h020, 16'h040, 16'h040, 16'h040, 16'h040, 16'h020, 16'h020, 16'h040, 16'h020, 16'h020, 16'h020, 16'h020, 16'h00, 16'h020, 16'h20e3, 16'h3164, 16'h2943, 16'h840, 16'h020, 16'h020, 16'h020, 16'h020, 16'h1081, 16'h213, 16'h3124, 16'h72ea, 16'h6247, 16'h6267, 16'h6267, 16'h6267, 16'h6267, 16'h6267, 16'h6267, 16'h6268, 16'h6288, 16'h6aa8, 16'h832a, 16'h9cd, 16'h5a67, 16'h3164, 16'h820, 16'h020, 16'h020, 16'h020, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h040, 16'h840, 16'h841, 16'h62a9, 16'hb512, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha470, 16'ha470, 16'ha46f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c4e, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9ce, 16'h9ce, 16'h9c2e, 16'h94e, 16'h94e, 16'h7b2b, 16'h3144, 16'h20c3, 16'h20c2, 16'h20c1, 16'h20c2, 16'h1061, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h732a, 16'h7b2a, 16'h7b4b, 16'h7b4b, 16'h7b6b, 16'h7b6b, 16'h836b, 16'h838b, 16'h838b, 16'h83ab, 16'h83ac, 16'h8bac, 16'h8bcc, 16'h8bcc, 16'h8bed, 16'h8bed, 16'h94d, 16'h94d, 16'h942e, 16'h9c2e, 16'h9c4e, 16'h944e, 16'h4a5, 16'h10a0, 16'h860, 16'h860, 16'h860, 16'h860, 16'h860, 16'h860, 16'h860, 16'h860, 16'h860, 16'h860, 16'h040, 16'h040, 16'h2923, 16'h5247, 16'h1081, 16'h860, 16'h840, 16'h020, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h020, 16'h020, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h020, 16'h040, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h18c2, 16'h3144, 16'h2943, 16'h840, 16'h020, 16'h020, 16'h020, 16'h020, 16'h18a2, 16'h2944, 16'h2923, 16'h73a, 16'h6248, 16'h6267, 16'h6267, 16'h6267, 16'h6267, 16'h6267, 16'h6267, 16'h6267, 16'h6a68, 16'h6aa8, 16'h832a, 16'h9cd, 16'h6267, 16'h3164, 16'h820, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h040, 16'h040, 16'h840, 16'h861, 16'h62a9, 16'hb512, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f2, 16'hb4d1, 16'hb4d1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb0, 16'hacb0, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4e, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h94e, 16'h94e, 16'h732b, 16'h3144, 16'h20e2, 16'h20e2, 16'h20c1, 16'h20c1, 16'h1081, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h732a, 16'h7b2a, 16'h7b4a, 16'h7b4b, 16'h7b6a, 16'h7b6b, 16'h836b, 16'h836b, 16'h838b, 16'h83ac, 16'h83ac, 16'h8bcc, 16'h8bcc, 16'h8bec, 16'h8bed, 16'h8bed, 16'h94d, 16'h942d, 16'h942e, 16'h9c4e, 16'h9c4e, 16'h9c4e, 16'h4a26, 16'h10a0, 16'h860, 16'h060, 16'h060, 16'h860, 16'h860, 16'h880, 16'h860, 16'h860, 16'h860, 16'h860, 16'h040, 16'h040, 16'h2923, 16'h5247, 16'h1081, 16'h860, 16'h020, 16'h020, 16'h040, 16'h040, 16'h020, 16'h040, 16'h040, 16'h040, 16'h020, 16'h020, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h820, 16'h861, 16'h1081, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h20c3, 16'h3985, 16'h293, 16'h73a, 16'h6268, 16'h6267, 16'h6267, 16'h5a67, 16'h6267, 16'h6267, 16'h6267, 16'h6267, 16'h6a87, 16'h6aa8, 16'h8329, 16'h9cd, 16'h6267, 16'h3164, 16'h820, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h040, 16'h040, 16'h840, 16'h860, 16'h62a9, 16'hb512, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c4e, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4e, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c4e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9ce, 16'h94e, 16'h7b4b, 16'h3144, 16'h20e2, 16'h20e2, 16'h20c1, 16'h20c1, 16'h1061, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h732a, 16'h7b2a, 16'h7b4a, 16'h7b4a, 16'h7b4b, 16'h7b6b, 16'h7b6b, 16'h838b, 16'h838b, 16'h83ac, 16'h83ab, 16'h83cc, 16'h8bcc, 16'h8bec, 16'h8bed, 16'h94d, 16'h94d, 16'h942e, 16'h942e, 16'h9c4e, 16'h9c4f, 16'h9c4e, 16'h4a26, 16'h10a1, 16'h060, 16'h060, 16'h860, 16'h860, 16'h860, 16'h860, 16'h860, 16'h060, 16'h060, 16'h060, 16'h040, 16'h020, 16'h2923, 16'h4a6, 16'h1081, 16'h840, 16'h020, 16'h840, 16'h040, 16'h040, 16'h020, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h040, 16'h020, 16'h020, 16'h293, 16'h41c6, 16'h294, 16'h732a, 16'h6267, 16'h5a67, 16'h6267, 16'h6267, 16'h6267, 16'h6267, 16'h6268, 16'h6267, 16'h6267, 16'h6aa8, 16'h8329, 16'h9cd, 16'h6267, 16'h3164, 16'h820, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h040, 16'h040, 16'h040, 16'h840, 16'h861, 16'h6aa9, 16'hb512, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb511, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha470, 16'ha470, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha44f, 16'h9c4f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c4f, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h94e, 16'h7b2b, 16'h3144, 16'h20e2, 16'h20e1, 16'h18c1, 16'h18c1, 16'h1080, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h732a, 16'h7b2a, 16'h7b2a, 16'h7b4a, 16'h7b4b, 16'h7b4b, 16'h836b, 16'h838b, 16'h838c, 16'h838c, 16'h83ab, 16'h83ac, 16'h8bcc, 16'h8bec, 16'h8bed, 16'h94d, 16'h942d, 16'h942e, 16'h9c4e, 16'h9c4e, 16'h9c6e, 16'h9c4e, 16'h5226, 16'h1081, 16'h060, 16'h060, 16'h860, 16'h860, 16'h880, 16'h880, 16'h860, 16'h860, 16'h060, 16'h060, 16'h040, 16'h040, 16'h3164, 16'h49e6, 16'h1081, 16'h840, 16'h820, 16'h840, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h040, 16'h020, 16'h3144, 16'h4a7, 16'h294, 16'h73a, 16'h6267, 16'h5a67, 16'h5a67, 16'h6267, 16'h6267, 16'h6267, 16'h5a67, 16'h6267, 16'h6267, 16'h6aa8, 16'h7b29, 16'h9cc, 16'h6267, 16'h3164, 16'h820, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h040, 16'h040, 16'h840, 16'h861, 16'h6aa9, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4e, 16'h9c4e, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c4f, 16'h9c4e, 16'h9c4e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9ce, 16'h7b2b, 16'h3144, 16'h20e2, 16'h20c2, 16'h20c1, 16'h20c1, 16'h1080, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h732a, 16'h7b2a, 16'h7b2a, 16'h7b4a, 16'h7b4b, 16'h7b4b, 16'h836b, 16'h838b, 16'h838b, 16'h838c, 16'h83ac, 16'h83ac, 16'h8bcc, 16'h8bcc, 16'h93ed, 16'h94d, 16'h94d, 16'h942e, 16'h9c2e, 16'h9c4e, 16'h9c6e, 16'h9c4e, 16'h5226, 16'h10a1, 16'h060, 16'h860, 16'h860, 16'h860, 16'h860, 16'h860, 16'h860, 16'h860, 16'h060, 16'h060, 16'h040, 16'h040, 16'h2944, 16'h41c5, 16'h1080, 16'h020, 16'h840, 16'h840, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h020, 16'h020, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h020, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h840, 16'h040, 16'h040, 16'h820, 16'h3164, 16'h49e6, 16'h294, 16'h7ba, 16'h6267, 16'h6267, 16'h6267, 16'h6267, 16'h6267, 16'h6267, 16'h6267, 16'h6267, 16'h6267, 16'h6aa8, 16'h7b29, 16'h9cc, 16'h6267, 16'h3164, 16'h820, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h040, 16'h040, 16'h040, 16'h840, 16'h1061, 16'h62a9, 16'hb512, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'ha490, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha46f, 16'ha46f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4e, 16'h9c4f, 16'h9c4f, 16'h9c2e, 16'h9c2e, 16'h9ce, 16'h7b4b, 16'h3144, 16'h20e2, 16'h20c2, 16'h20c1, 16'h18c1, 16'h1080, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h7329, 16'h7b2a, 16'h7b4a, 16'h7b4b, 16'h7b4b, 16'h7b6b, 16'h836b, 16'h838b, 16'h838c, 16'h838c, 16'h83ac, 16'h83ac, 16'h8bcc, 16'h8bcc, 16'h8bec, 16'h94d, 16'h94d, 16'h942e, 16'h9c2e, 16'h9c4e, 16'h9c4e, 16'h9c4e, 16'h5246, 16'h10a0, 16'h860, 16'h880, 16'h880, 16'h880, 16'h860, 16'h860, 16'h860, 16'h860, 16'h860, 16'h860, 16'h040, 16'h040, 16'h213, 16'h3184, 16'h860, 16'h861, 16'h1081, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h020, 16'h020, 16'h040, 16'h040, 16'h040, 16'h020, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h840, 16'h840, 16'h860, 16'h1081, 16'h1081, 16'h1061, 16'h1061, 16'h3165, 16'h41c5, 16'h20e3, 16'h73a, 16'h6267, 16'h6267, 16'h6267, 16'h6267, 16'h6267, 16'h6267, 16'h6267, 16'h6267, 16'h6267, 16'h6a88, 16'h8329, 16'h9cc, 16'h6267, 16'h3164, 16'h820, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h820, 16'h020, 16'h020, 16'h040, 16'h040, 16'h040, 16'h840, 16'h1061, 16'h6aa9, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'ha490, 16'hac90, 16'hac90, 16'hac90, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha46f, 16'ha470, 16'ha470, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9ce, 16'h7b4b, 16'h3164, 16'h20e2, 16'h20e2, 16'h20c1, 16'h20c2, 16'h1081, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h739, 16'h732a, 16'h7b4a, 16'h7b4a, 16'h7b4b, 16'h7b6b, 16'h7b6b, 16'h838b, 16'h838b, 16'h838c, 16'h83ac, 16'h83ac, 16'h8bcc, 16'h8bcc, 16'h8bed, 16'h93ed, 16'h94d, 16'h942d, 16'h9c2e, 16'h9c4e, 16'h9c4f, 16'h9c4e, 16'h4a26, 16'h1081, 16'h861, 16'h880, 16'h880, 16'h880, 16'h880, 16'h880, 16'h860, 16'h860, 16'h860, 16'h860, 16'h860, 16'h860, 16'h10c1, 16'h212, 16'h860, 16'h860, 16'h860, 16'h840, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h020, 16'h040, 16'h040, 16'h040, 16'h020, 16'h020, 16'h040, 16'h020, 16'h040, 16'h020, 16'h040, 16'h020, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h840, 16'h861, 16'h1081, 16'h18a2, 16'h18a1, 16'h18a2, 16'h3985, 16'h41e6, 16'h3124, 16'h72ea, 16'h6267, 16'h6267, 16'h6267, 16'h6267, 16'h6267, 16'h6267, 16'h6267, 16'h6267, 16'h6a68, 16'h6a88, 16'h839, 16'h9cc, 16'h6267, 16'h3964, 16'h820, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h040, 16'h040, 16'h040, 16'h840, 16'h1061, 16'h6aa9, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd0, 16'hacd0, 16'hacb0, 16'hacb0, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'hac90, 16'hac90, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha470, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha470, 16'ha450, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c2e, 16'h7b4b, 16'h3144, 16'h20e2, 16'h20c2, 16'h20c1, 16'h20c1, 16'h1081, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h7329, 16'h732a, 16'h7b2a, 16'h7b4a, 16'h7b4a, 16'h7b4b, 16'h7b6b, 16'h836b, 16'h838b, 16'h838c, 16'h83ac, 16'h83ac, 16'h8bcc, 16'h8bcc, 16'h8bed, 16'h93ed, 16'h94d, 16'h942e, 16'h9c2e, 16'h9c4e, 16'h9c4e, 16'h9c4e, 16'h4a26, 16'h1081, 16'h860, 16'h860, 16'h860, 16'h880, 16'h880, 16'h860, 16'h860, 16'h860, 16'h860, 16'h860, 16'h860, 16'h860, 16'h860, 16'h060, 16'h060, 16'h10a1, 16'h41c5, 16'h41c5, 16'h3144, 16'h20e3, 16'h18a2, 16'h1081, 16'h860, 16'h040, 16'h040, 16'h020, 16'h040, 16'h020, 16'h020, 16'h040, 16'h040, 16'h040, 16'h020, 16'h020, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h860, 16'h860, 16'h1881, 16'h1882, 16'h20e3, 16'h3144, 16'h2924, 16'h214, 16'h72ea, 16'h6248, 16'h6248, 16'h6267, 16'h6267, 16'h6267, 16'h6267, 16'h6267, 16'h6267, 16'h6267, 16'h6a88, 16'h7ba, 16'h9cc, 16'h6267, 16'h3964, 16'h820, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h040, 16'h040, 16'h040, 16'h040, 16'h840, 16'h861, 16'h62a9, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd0, 16'hacd0, 16'hacb0, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'hac90, 16'hac90, 16'hac90, 16'hac90, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha46f, 16'ha46f, 16'ha470, 16'ha470, 16'ha46f, 16'ha46f, 16'ha470, 16'ha46f, 16'ha470, 16'ha46f, 16'ha450, 16'ha44f, 16'ha44f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'h9c4f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c2e, 16'h7b4b, 16'h3164, 16'h20e2, 16'h20e2, 16'h20c1, 16'h20c1, 16'h1080, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h7329, 16'h732a, 16'h7b2a, 16'h7b4a, 16'h7b4b, 16'h7b6b, 16'h7b6b, 16'h838b, 16'h838c, 16'h838b, 16'h83ab, 16'h83ac, 16'h8bcc, 16'h8bec, 16'h8bed, 16'h93ed, 16'h94d, 16'h94e, 16'h942e, 16'h9c4e, 16'h9c4f, 16'h9c4e, 16'h73a, 16'h49e6, 16'h39a5, 16'h2964, 16'h213, 16'h18e2, 16'h10a1, 16'h881, 16'h880, 16'h860, 16'h860, 16'h860, 16'h860, 16'h860, 16'h860, 16'h060, 16'h060, 16'h10a1, 16'h72e9, 16'h838b, 16'h836b, 16'h7b2a, 16'h73a, 16'h6ae9, 16'h49e5, 16'h881, 16'h860, 16'h10a2, 16'h1081, 16'h840, 16'h040, 16'h840, 16'h040, 16'h020, 16'h020, 16'h020, 16'h020, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h860, 16'h1081, 16'h1882, 16'h3165, 16'h2926, 16'h20e6, 16'h2926, 16'h73b, 16'h5a47, 16'h6248, 16'h6247, 16'h6267, 16'h5a67, 16'h6267, 16'h6247, 16'h6267, 16'h6267, 16'h6aa8, 16'h7b9, 16'h94c, 16'h5a67, 16'h3964, 16'h820, 16'h020, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h040, 16'h040, 16'h840, 16'h840, 16'h840, 16'h1061, 16'h62a9, 16'hb512, 16'hbd32, 16'hbd32, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha46f, 16'ha46f, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha450, 16'ha470, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c2e, 16'h7b4b, 16'h3144, 16'h20e2, 16'h20c2, 16'h20c2, 16'h20c1, 16'h1080, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h73a, 16'h732a, 16'h732a, 16'h7b4a, 16'h7b4b, 16'h7b4b, 16'h7b6b, 16'h838b, 16'h838b, 16'h838b, 16'h83ac, 16'h83ac, 16'h8bcc, 16'h8bec, 16'h8bec, 16'h94d, 16'h94d, 16'h942d, 16'h942e, 16'h944e, 16'h9c4e, 16'h9c4f, 16'h9c4f, 16'h9c4e, 16'h9c4e, 16'h9c4e, 16'h94e, 16'h8bed, 16'h83ac, 16'h7b6b, 16'h6ba, 16'h62c9, 16'h5248, 16'h39c5, 16'h213, 16'h20e2, 16'h18c2, 16'h18a1, 16'h881, 16'h18a1, 16'h72e9, 16'h8bab, 16'h8bab, 16'h8b8c, 16'h8bac, 16'h93ec, 16'h6ac8, 16'h1061, 16'h1081, 16'h41c6, 16'h3164, 16'h20e3, 16'h18c2, 16'h18a2, 16'h10a1, 16'h1081, 16'h861, 16'h861, 16'h840, 16'h840, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h860, 16'h861, 16'h293, 16'h5a8b, 16'h214a, 16'h199, 16'h3168, 16'h7ba, 16'h6247, 16'h6248, 16'h6247, 16'h6247, 16'h5a47, 16'h6247, 16'h6247, 16'h6267, 16'h6267, 16'h6aa8, 16'h7ba, 16'h9cc, 16'h5a67, 16'h3164, 16'h820, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h040, 16'h040, 16'h840, 16'h840, 16'h840, 16'h1061, 16'h6aa9, 16'hb512, 16'hbd32, 16'hbd32, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd0, 16'hacd0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha470, 16'ha46f, 16'ha46f, 16'ha470, 16'ha470, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha46f, 16'ha46f, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha46f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c2e, 16'h7b4b, 16'h3144, 16'h20e2, 16'h20c2, 16'h20c2, 16'h20c2, 16'h1081, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h73a, 16'h732a, 16'h7b4a, 16'h7b4a, 16'h7b4b, 16'h7b6b, 16'h7b6b, 16'h838b, 16'h838b, 16'h838b, 16'h83ac, 16'h83ac, 16'h83cc, 16'h8bcc, 16'h8bed, 16'h94d, 16'h94d, 16'h942d, 16'h942e, 16'h944e, 16'h9c4e, 16'h9c4f, 16'h9c6f, 16'h9c6f, 16'ha46f, 16'ha48f, 16'ha4af, 16'ha4b0, 16'ha4b0, 16'hacb0, 16'hacd0, 16'hacb0, 16'hacb0, 16'h8bec, 16'h6aa8, 16'h6287, 16'h5a67, 16'h5a67, 16'h41c5, 16'h3123, 16'h6aa8, 16'h7b4a, 16'h836b, 16'h8bab, 16'h93ac, 16'h94c, 16'h6ac8, 16'h1081, 16'h1881, 16'h4a7, 16'h3985, 16'h2924, 16'h213, 16'h213, 16'h213, 16'h213, 16'h20e3, 16'h20e3, 16'h18c3, 16'h18c2, 16'h10a2, 16'h1081, 16'h1061, 16'h861, 16'h840, 16'h861, 16'h861, 16'h040, 16'h040, 16'h040, 16'h040, 16'h841, 16'h214, 16'h42c, 16'h216b, 16'h296b, 16'h2928, 16'h7ae9, 16'h6a68, 16'h5a47, 16'h5a67, 16'h6247, 16'h5a47, 16'h6267, 16'h6267, 16'h6267, 16'h6a68, 16'h6aa8, 16'h7b9, 16'h9bec, 16'h5a67, 16'h3164, 16'h020, 16'h020, 16'h840, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h040, 16'h040, 16'h840, 16'h840, 16'h840, 16'h1061, 16'h6aa9, 16'hbd12, 16'hbd32, 16'hbd32, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f2, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha46f, 16'ha470, 16'ha46f, 16'ha470, 16'ha470, 16'ha450, 16'ha44f, 16'ha44f, 16'h9c2f, 16'h7b4b, 16'h3144, 16'h20e2, 16'h20c2, 16'h20c2, 16'h20c2, 16'h1081, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h732a, 16'h7b2a, 16'h7b4a, 16'h7b4a, 16'h7b4a, 16'h7b6b, 16'h7b8b, 16'h838b, 16'h838b, 16'h838c, 16'h83ac, 16'h83ac, 16'h8bcc, 16'h8bcc, 16'h8bed, 16'h93ed, 16'h94d, 16'h94d, 16'h942e, 16'h944e, 16'h9c4e, 16'h9c4e, 16'h9c4f, 16'h9c6f, 16'h9c6f, 16'h9c6f, 16'ha48f, 16'ha48f, 16'ha4af, 16'ha4af, 16'h9c6e, 16'h8bed, 16'h7b8b, 16'h62c8, 16'h49e6, 16'h41c5, 16'h3985, 16'h3964, 16'h3164, 16'h3124, 16'h3964, 16'h3984, 16'h41c5, 16'h6288, 16'h8bac, 16'h94c, 16'h6ae8, 16'h1081, 16'h18a2, 16'h49e6, 16'h3164, 16'h2923, 16'h213, 16'h213, 16'h213, 16'h213, 16'h213, 16'h213, 16'h213, 16'h213, 16'h213, 16'h213, 16'h213, 16'h20e3, 16'h18c2, 16'h18c3, 16'h18c2, 16'h10a2, 16'h10a2, 16'h1081, 16'h861, 16'h862, 16'h10c6, 16'h212b, 16'h298b, 16'h39a9, 16'h3126, 16'h839, 16'h6a88, 16'h5a47, 16'h5a47, 16'h5a47, 16'h5a47, 16'h6247, 16'h5a47, 16'h6267, 16'h6268, 16'h6aa8, 16'h7b9, 16'h93ec, 16'h6267, 16'h3164, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h840, 16'h1061, 16'h6aa9, 16'hbd12, 16'hbd32, 16'hbd32, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha44f, 16'h9c4f, 16'h7b6b, 16'h3164, 16'h20e2, 16'h20c2, 16'h20c2, 16'h20c2, 16'h1081, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h732a, 16'h7b4a, 16'h7b4a, 16'h7b4b, 16'h7b4b, 16'h7b6b, 16'h836b, 16'h838b, 16'h838c, 16'h838c, 16'h83ac, 16'h83ac, 16'h8bcc, 16'h8bcd, 16'h8bed, 16'h8cd, 16'h94d, 16'h942d, 16'h942d, 16'h942e, 16'h9c4e, 16'h9c4e, 16'h9c6e, 16'h9c6f, 16'h9c6f, 16'h9c6f, 16'h9c6f, 16'h9c4e, 16'h942d, 16'h7b4a, 16'h5a67, 16'h41c5, 16'h3164, 16'h3144, 16'h2924, 16'h293, 16'h293, 16'h28e3, 16'h20e3, 16'h20e3, 16'h20e3, 16'h213, 16'h20e3, 16'h2923, 16'h6287, 16'h94c, 16'h6ae8, 16'h1081, 16'h18a2, 16'h41e6, 16'h3165, 16'h2924, 16'h293, 16'h293, 16'h294, 16'h214, 16'h293, 16'h2923, 16'h293, 16'h213, 16'h213, 16'h2923, 16'h2923, 16'h2924, 16'h293, 16'h293, 16'h2924, 16'h2924, 16'h294, 16'h2924, 16'h214, 16'h18e5, 16'h192a, 16'h216c, 16'h39ca, 16'h4a28, 16'h49c5, 16'h8b48, 16'h6a87, 16'h5a47, 16'h6247, 16'h6247, 16'h5a47, 16'h5a47, 16'h5a47, 16'h6247, 16'h6267, 16'h6aa8, 16'h7b9, 16'h93ec, 16'h6267, 16'h3164, 16'h820, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h040, 16'h040, 16'h040, 16'h040, 16'h840, 16'h840, 16'h1061, 16'h6aa9, 16'hbd12, 16'hbd32, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'ha490, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha48f, 16'ha48f, 16'ha490, 16'ha46f, 16'ha46f, 16'ha470, 16'ha470, 16'ha46f, 16'ha46f, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha46f, 16'ha46f, 16'h9c4f, 16'h836c, 16'h3164, 16'h20e2, 16'h20c2, 16'h20c1, 16'h20c1, 16'h1081, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h732a, 16'h7b4a, 16'h7b4a, 16'h7b4a, 16'h7b6a, 16'h7b6b, 16'h836b, 16'h838c, 16'h838c, 16'h83ac, 16'h83ac, 16'h83ac, 16'h8bcc, 16'h8bcc, 16'h8bed, 16'h8bed, 16'h94d, 16'h942d, 16'h942e, 16'h942e, 16'h9c4e, 16'h9c4e, 16'h9c4e, 16'h9c6f, 16'h9c6f, 16'h9c6f, 16'h9c6e, 16'h838b, 16'h5a87, 16'h4184, 16'h3144, 16'h2924, 16'h2923, 16'h293, 16'h213, 16'h293, 16'h28e3, 16'h20e3, 16'h20c3, 16'h20e3, 16'h20e3, 16'h20e3, 16'h20e3, 16'h20c2, 16'h3984, 16'h93cc, 16'h6ae8, 16'h1081, 16'h18c2, 16'h41e6, 16'h3965, 16'h2924, 16'h2923, 16'h293, 16'h293, 16'h294, 16'h2923, 16'h2923, 16'h293, 16'h293, 16'h213, 16'h293, 16'h293, 16'h293, 16'h294, 16'h2924, 16'h2924, 16'h2924, 16'h2925, 16'h62ca, 16'h62aa, 16'h2947, 16'h212a, 16'h294a, 16'h4aa, 16'h6aaa, 16'h7ba, 16'h9389, 16'h5a25, 16'h526, 16'h5a26, 16'h5a26, 16'h5a46, 16'h5a46, 16'h5a47, 16'h5a47, 16'h6267, 16'h6a88, 16'h7b9, 16'h93ec, 16'h5a67, 16'h3964, 16'h840, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h040, 16'h040, 16'h040, 16'h840, 16'h840, 16'h840, 16'h1061, 16'h6aa9, 16'hbd12, 16'hbd32, 16'hbd32, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'hac90, 16'ha490, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha48f, 16'ha48f, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha46f, 16'ha44f, 16'h836c, 16'h3164, 16'h20e3, 16'h20c2, 16'h20c2, 16'h20c2, 16'h1081, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h7b2a, 16'h7b4a, 16'h7b6a, 16'h7b6b, 16'h7b6b, 16'h7b6b, 16'h836b, 16'h838c, 16'h838b, 16'h83ab, 16'h83ac, 16'h83ad, 16'h8bcc, 16'h8bec, 16'h8bed, 16'h8cd, 16'h94d, 16'h942d, 16'h942e, 16'h942e, 16'h9c2e, 16'h9c4e, 16'h9c4e, 16'h9c6e, 16'h9c6f, 16'h9c6f, 16'h8bcc, 16'h5a68, 16'h3985, 16'h3123, 16'h293, 16'h293, 16'h213, 16'h293, 16'h20e3, 16'h20e3, 16'h20e3, 16'h20e2, 16'h20c3, 16'h20c3, 16'h20c2, 16'h20e2, 16'h20c2, 16'h18a2, 16'h28e3, 16'h838b, 16'h6ae8, 16'h1081, 16'h20e3, 16'h41c5, 16'h3964, 16'h2924, 16'h2923, 16'h293, 16'h293, 16'h293, 16'h2923, 16'h2924, 16'h2924, 16'h2924, 16'h294, 16'h293, 16'h293, 16'h293, 16'h2923, 16'h2924, 16'h2924, 16'h2924, 16'h3986, 16'h942f, 16'h7b6d, 16'h2127, 16'h18e9, 16'h294a, 16'h41ea, 16'h628a, 16'h93cd, 16'h72c8, 16'h51e4, 16'h51c4, 16'h49c4, 16'h51c3, 16'h51e3, 16'h5a4, 16'h5a24, 16'h5a25, 16'h6245, 16'h6a66, 16'h7b8, 16'h93ec, 16'h5a67, 16'h3984, 16'h18c2, 16'h20c2, 16'h212, 16'h212, 16'h20c2, 16'h18a1, 16'h1081, 16'h861, 16'h840, 16'h840, 16'h820, 16'h840, 16'h840, 16'h020, 16'h840, 16'h840, 16'h040, 16'h840, 16'h840, 16'h840, 16'h1061, 16'h6aaa, 16'hbd12, 16'hbd12, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'hac90, 16'hac90, 16'ha490, 16'hac90, 16'ha490, 16'hac90, 16'hac90, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha48f, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha490, 16'ha490, 16'ha470, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha490, 16'ha470, 16'ha470, 16'ha46f, 16'ha44f, 16'h7b6c, 16'h3164, 16'h20e2, 16'h20c2, 16'h20c2, 16'h20c1, 16'h1081, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h7b4a, 16'h7b6a, 16'h7b6a, 16'h7b6b, 16'h836b, 16'h838b, 16'h838c, 16'h838c, 16'h83ac, 16'h83ac, 16'h83ac, 16'h8bcc, 16'h8bcc, 16'h8bed, 16'h8bed, 16'h94d, 16'h94d, 16'h942e, 16'h942e, 16'h9c2e, 16'h9c4e, 16'h9c4e, 16'h9c6f, 16'h9c6f, 16'h9c6f, 16'h94d, 16'h62c9, 16'h41c5, 16'h3144, 16'h293, 16'h213, 16'h20e3, 16'h20e3, 16'h20e2, 16'h20e3, 16'h20e3, 16'h20c3, 16'h20c3, 16'h20c2, 16'h20c2, 16'h20c2, 16'h20a2, 16'h18a2, 16'h18a1, 16'h1881, 16'h5a47, 16'h5a67, 16'h18c2, 16'h293, 16'h3144, 16'h3144, 16'h2923, 16'h293, 16'h294, 16'h294, 16'h293, 16'h294, 16'h2924, 16'h2924, 16'h2924, 16'h293, 16'h2923, 16'h2923, 16'h2924, 16'h2923, 16'h2924, 16'h2944, 16'h3144, 16'h4a8, 16'ha4b1, 16'h732c, 16'h2927, 16'h212a, 16'h2129, 16'h18c7, 16'h62ab, 16'h8b8c, 16'h5a27, 16'h526, 16'h51e5, 16'h49c5, 16'h49a4, 16'h49a4, 16'h49c4, 16'h51e4, 16'h51e4, 16'h5a4, 16'h6a45, 16'h7ac7, 16'h8baa, 16'h5a66, 16'h3984, 16'h18c1, 16'h212, 16'h3983, 16'h41c4, 16'h49e5, 16'h49e5, 16'h41c4, 16'h41a4, 16'h3984, 16'h3163, 16'h2923, 16'h20e2, 16'h20c2, 16'h1881, 16'h1081, 16'h861, 16'h840, 16'h840, 16'h840, 16'h840, 16'h1061, 16'h6aa9, 16'hbd12, 16'hbd12, 16'hbd32, 16'hbd32, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f2, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacd0, 16'hacb0, 16'hacb0, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hacb0, 16'hac90, 16'hac90, 16'ha490, 16'hac90, 16'ha490, 16'hac90, 16'hac90, 16'hac90, 16'hac90, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha450, 16'h836c, 16'h3164, 16'h20e2, 16'h20e2, 16'h20c2, 16'h20c2, 16'h1081, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h7b4a, 16'h7b6a, 16'h7b6b, 16'h7b6b, 16'h836b, 16'h838c, 16'h838c, 16'h838c, 16'h83ac, 16'h83ac, 16'h83ac, 16'h8bcc, 16'h8bec, 16'h8bed, 16'h94d, 16'h94d, 16'h942d, 16'h942e, 16'h942e, 16'h9c4e, 16'h9c4f, 16'h9c4f, 16'h9c6f, 16'h9c6f, 16'h9c6e, 16'h7b4a, 16'h49e6, 16'h3965, 16'h2943, 16'h293, 16'h293, 16'h213, 16'h20e3, 16'h20e3, 16'h20e3, 16'h20e3, 16'h20c3, 16'h20c3, 16'h20c2, 16'h18a2, 16'h18a1, 16'h1881, 16'h1081, 16'h881, 16'h1060, 16'h20c2, 16'h3123, 16'h2923, 16'h2923, 16'h3144, 16'h3144, 16'h2923, 16'h2923, 16'h294, 16'h294, 16'h2923, 16'h294, 16'h294, 16'h2924, 16'h2923, 16'h2924, 16'h2923, 16'h2923, 16'h2924, 16'h2923, 16'h2923, 16'h2944, 16'h3144, 16'h4a28, 16'h8bee, 16'h5228, 16'h2928, 16'h296a, 16'h18e8, 16'h18c7, 16'h732c, 16'h6aa9, 16'h5227, 16'h5a27, 16'h5227, 16'h526, 16'h49e5, 16'h49c5, 16'h49c5, 16'h49c5, 16'h49e5, 16'h5a27, 16'h6aa8, 16'h8b8a, 16'h739, 16'h41c5, 16'h20e2, 16'h820, 16'h840, 16'h1061, 16'h18a1, 16'h18c2, 16'h212, 16'h2943, 16'h3183, 16'h39a4, 16'h41c4, 16'h49e5, 16'h4a5, 16'h49e5, 16'h49e5, 16'h41c5, 16'h39a4, 16'h3984, 16'h3143, 16'h2923, 16'h20e2, 16'h20c2, 16'h6aca, 16'hbd12, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacd1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'hac90, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'hac90, 16'hac90, 16'hacb0, 16'hac90, 16'ha490, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'h838c, 16'h3164, 16'h20e2, 16'h20e2, 16'h20c2, 16'h18c2, 16'h1081, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h7b4a, 16'h836b, 16'h836b, 16'h836b, 16'h838b, 16'h838c, 16'h838c, 16'h83ac, 16'h83ac, 16'h83ac, 16'h8bcd, 16'h8bcd, 16'h8bed, 16'h8cd, 16'h94d, 16'h942d, 16'h942d, 16'h942e, 16'h9c4e, 16'h9c4e, 16'h9c4f, 16'h9c6f, 16'h9c6f, 16'h9c6f, 16'h9c4e, 16'h62c9, 16'h41c5, 16'h3164, 16'h3144, 16'h2923, 16'h293, 16'h213, 16'h213, 16'h213, 16'h20e3, 16'h20e3, 16'h20e2, 16'h20c2, 16'h18a2, 16'h18a1, 16'h1081, 16'h861, 16'h860, 16'h860, 16'h860, 16'h1060, 16'h1881, 16'h18c1, 16'h20e2, 16'h3144, 16'h2944, 16'h2923, 16'h2923, 16'h2923, 16'h2924, 16'h2924, 16'h294, 16'h294, 16'h294, 16'h2923, 16'h2924, 16'h2923, 16'h2924, 16'h2924, 16'h2923, 16'h2924, 16'h2944, 16'h2944, 16'h3144, 16'h41c6, 16'h3165, 16'h2947, 16'h216, 16'h18a4, 16'h20e5, 16'h5a68, 16'h5a47, 16'h5a46, 16'h5a46, 16'h5a47, 16'h5a27, 16'h5226, 16'h526, 16'h49c5, 16'h49c5, 16'h49e6, 16'h5a47, 16'h832a, 16'h836a, 16'h524, 16'h2922, 16'h840, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h820, 16'h840, 16'h860, 16'h1061, 16'h18a1, 16'h18c1, 16'h212, 16'h2943, 16'h3163, 16'h39a4, 16'h41c4, 16'h49e5, 16'h49e5, 16'h4a5, 16'h526, 16'h836c, 16'hbd12, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'hac90, 16'hac90, 16'hac90, 16'hac90, 16'hac90, 16'hacb0, 16'hacb0, 16'hac90, 16'hacb0, 16'hac90, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'h838c, 16'h3965, 16'h20e3, 16'h20c2, 16'h20c2, 16'h18c2, 16'h1081, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h7b4a, 16'h7b6a, 16'h838b, 16'h838b, 16'h838b, 16'h838c, 16'h83ac, 16'h83ac, 16'h83ac, 16'h8bcc, 16'h8bcc, 16'h8bed, 16'h8bed, 16'h94d, 16'h94d, 16'h942d, 16'h942e, 16'h9c4e, 16'h9c4e, 16'h9c6f, 16'h9c6f, 16'h9c6f, 16'ha48f, 16'ha48f, 16'h9c4f, 16'h62a8, 16'h41c5, 16'h3164, 16'h2924, 16'h294, 16'h293, 16'h293, 16'h213, 16'h20e3, 16'h20e3, 16'h20e2, 16'h20e2, 16'h18c2, 16'h18a2, 16'h1081, 16'h860, 16'h860, 16'h860, 16'h860, 16'h860, 16'h840, 16'h840, 16'h840, 16'h20c2, 16'h3964, 16'h3144, 16'h2923, 16'h2923, 16'h2924, 16'h2924, 16'h2924, 16'h294, 16'h294, 16'h2924, 16'h2923, 16'h2924, 16'h2924, 16'h2923, 16'h2923, 16'h2923, 16'h2923, 16'h2924, 16'h3144, 16'h2944, 16'h2924, 16'h20e2, 16'h1081, 16'h841, 16'h841, 16'h1061, 16'h20e2, 16'h4185, 16'h5227, 16'h5a47, 16'h5a47, 16'h5a47, 16'h5a47, 16'h5226, 16'h5226, 16'h5226, 16'h5a47, 16'h6ac9, 16'h8bab, 16'h5a66, 16'h3163, 16'h1081, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h820, 16'h820, 16'h840, 16'h840, 16'h1080, 16'h18a1, 16'h18c1, 16'h28e2, 16'h3123, 16'h7b2a, 16'hbd12, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hbd32, 16'hbd12, 16'hbd12, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f2, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'ha44f, 16'h9c4f, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'hac90, 16'hac90, 16'hac90, 16'hac90, 16'hac90, 16'hac90, 16'hac90, 16'hac90, 16'hac90, 16'hac90, 16'hacb0, 16'hac90, 16'hacb0, 16'hacb0, 16'hacb0, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'h838c, 16'h3165, 16'h20e3, 16'h20e2, 16'h20c1, 16'h18c2, 16'h1061, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h6ae9, 16'h6b9, 16'h739, 16'h7329, 16'h732a, 16'h7b4a, 16'h7b6b, 16'h838b, 16'h83ac, 16'h83cc, 16'h8bcd, 16'h8bed, 16'h94d, 16'h94d, 16'h942d, 16'h944d, 16'h9c4e, 16'h9c4e, 16'h9c6e, 16'h9c4e, 16'h9c6f, 16'h9c8f, 16'ha48f, 16'ha48f, 16'h9c6e, 16'h62a8, 16'h39a5, 16'h3164, 16'h2924, 16'h293, 16'h20e3, 16'h20e3, 16'h20e3, 16'h20e3, 16'h20e3, 16'h20e3, 16'h20c3, 16'h20c3, 16'h18a2, 16'h860, 16'h060, 16'h060, 16'h060, 16'h860, 16'h840, 16'h020, 16'h020, 16'h020, 16'h18a2, 16'h3985, 16'h3144, 16'h2924, 16'h2924, 16'h2924, 16'h2923, 16'h2924, 16'h2924, 16'h2924, 16'h2924, 16'h2923, 16'h2923, 16'h2923, 16'h2923, 16'h2123, 16'h2923, 16'h2923, 16'h2944, 16'h3144, 16'h2944, 16'h2944, 16'h213, 16'h840, 16'h020, 16'h861, 16'h840, 16'h840, 16'h1061, 16'h2923, 16'h49c5, 16'h526, 16'h5227, 16'h5227, 16'h5227, 16'h5a47, 16'h6267, 16'h72c9, 16'h8bac, 16'h6ac8, 16'h3142, 16'h18a1, 16'h020, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h040, 16'h040, 16'h840, 16'h840, 16'h1041, 16'h6aa9, 16'hbd12, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hbd32, 16'hbd32, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f2, 16'hb4f1, 16'ha490, 16'h732b, 16'h527, 16'h49e6, 16'h7b4b, 16'hacd0, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'hac90, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hacb0, 16'hacb0, 16'hacb0, 16'ha490, 16'hacb0, 16'hac90, 16'ha470, 16'h838c, 16'h3165, 16'h20e3, 16'h20c2, 16'h20c2, 16'h20c2, 16'h1061, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h7b6b, 16'h838b, 16'h838b, 16'h7b6b, 16'h7b6a, 16'h7b4a, 16'h7b4a, 16'h734a, 16'h732a, 16'h7b4a, 16'h7b4a, 16'h7b6b, 16'h83ac, 16'h8bcc, 16'h8bed, 16'h942d, 16'h942e, 16'h9c4f, 16'h942e, 16'h5a88, 16'h5247, 16'h6b9, 16'h7b8b, 16'h8bed, 16'h942d, 16'h62a9, 16'h3985, 16'h3164, 16'h2924, 16'h213, 16'h20e3, 16'h20c2, 16'h20c2, 16'h20e2, 16'h20e2, 16'h20e3, 16'h20c3, 16'h20c3, 16'h20c2, 16'h1081, 16'h860, 16'h060, 16'h060, 16'h840, 16'h040, 16'h020, 16'h040, 16'h840, 16'h18a2, 16'h3985, 16'h3144, 16'h2923, 16'h2923, 16'h293, 16'h293, 16'h294, 16'h2923, 16'h293, 16'h294, 16'h2923, 16'h2924, 16'h2923, 16'h2923, 16'h2123, 16'h213, 16'h293, 16'h2923, 16'h2924, 16'h2924, 16'h3164, 16'h2924, 16'h840, 16'h1081, 16'h41e6, 16'h18a2, 16'h040, 16'h020, 16'h840, 16'h1081, 16'h20c2, 16'h294, 16'h3124, 16'h49e6, 16'h6288, 16'h6aa9, 16'h8b8b, 16'h838b, 16'h41a4, 16'h18c1, 16'h820, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h040, 16'h040, 16'h840, 16'h1061, 16'h6aaa, 16'hbd12, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb512, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hacb1, 16'h6aea, 16'h3165, 16'h3165, 16'h2924, 16'h41a6, 16'h9c2e, 16'hacd1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb1, 16'hacb0, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'hac90, 16'ha490, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'ha470, 16'h838d, 16'h3164, 16'h20e2, 16'h20c2, 16'h20c1, 16'h18c2, 16'h1081, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h838b, 16'h83ab, 16'h8bcc, 16'h8bcc, 16'h8bcc, 16'h8bcc, 16'h8bcc, 16'h8bec, 16'h8bec, 16'h8bcc, 16'h8bcc, 16'h8bcc, 16'h8bcc, 16'h8bcd, 16'h8bcc, 16'h8bcc, 16'h8bcd, 16'h8bcd, 16'h83ac, 16'h3164, 16'h1081, 16'h18c1, 16'h20e2, 16'h2923, 16'h3984, 16'h49e6, 16'h3985, 16'h3144, 16'h2923, 16'h20e3, 16'h20c2, 16'h20c2, 16'h20c2, 16'h20c2, 16'h20c2, 16'h20c2, 16'h20c3, 16'h20c2, 16'h20c2, 16'h18a1, 16'h1060, 16'h840, 16'h840, 16'h840, 16'h040, 16'h040, 16'h860, 16'h880, 16'h18a2, 16'h3985, 16'h3144, 16'h2923, 16'h2123, 16'h293, 16'h214, 16'h294, 16'h2923, 16'h293, 16'h293, 16'h214, 16'h293, 16'h2123, 16'h293, 16'h2923, 16'h293, 16'h293, 16'h2924, 16'h2924, 16'h2924, 16'h2924, 16'h1061, 16'h020, 16'h1081, 16'h41a4, 16'h1061, 16'h1082, 16'h841, 16'h020, 16'h020, 16'h840, 16'h861, 16'h18a3, 16'h4a6, 16'h73a, 16'h5226, 16'h5226, 16'h41c5, 16'h212, 16'h1881, 16'h840, 16'h840, 16'h820, 16'h020, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h040, 16'h040, 16'h040, 16'h861, 16'h6aa9, 16'hbd32, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hbd32, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f2, 16'hb4d1, 16'h7b4c, 16'h3165, 16'h2924, 16'h2924, 16'h2124, 16'h214, 16'h7b6c, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hac90, 16'ha470, 16'h838d, 16'h3164, 16'h20e2, 16'h20c2, 16'h20c2, 16'h18c2, 16'h1061, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h838b, 16'h8bab, 16'h8bcc, 16'h8bcc, 16'h8bcc, 16'h8bcc, 16'h8bed, 16'h8bed, 16'h8bed, 16'h94d, 16'h94d, 16'h942d, 16'h942d, 16'h944e, 16'h9c4e, 16'h9c6f, 16'h9c6f, 16'h9c8f, 16'h942e, 16'h3984, 16'h881, 16'h881, 16'h1080, 16'h1081, 16'h1881, 16'h3985, 16'h3985, 16'h3164, 16'h2923, 16'h20e2, 16'h18c2, 16'h18c2, 16'h18c2, 16'h20c2, 16'h18c2, 16'h20c2, 16'h18c2, 16'h20c2, 16'h20c2, 16'h20a2, 16'h18a2, 16'h1081, 16'h840, 16'h840, 16'h860, 16'h881, 16'h10a1, 16'h18c1, 16'h212, 16'h39a5, 16'h3144, 16'h2923, 16'h2923, 16'h2923, 16'h2924, 16'h294, 16'h2923, 16'h2924, 16'h294, 16'h2924, 16'h2924, 16'h2923, 16'h294, 16'h2923, 16'h293, 16'h213, 16'h294, 16'h2944, 16'h2944, 16'h213, 16'h861, 16'h020, 16'h1060, 16'h4142, 16'h4184, 16'h296, 16'h1085, 16'h843, 16'h041, 16'h020, 16'h020, 16'h840, 16'h1061, 16'h20c2, 16'h20c1, 16'h20c1, 16'h20c2, 16'h20e2, 16'h20e1, 16'h20c1, 16'h20c1, 16'h20c2, 16'h18c2, 16'h18a2, 16'h10a1, 16'h1081, 16'h1061, 16'h841, 16'h840, 16'h820, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h040, 16'h040, 16'h040, 16'h841, 16'h6aa9, 16'hbd32, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'h9c4f, 16'h49e7, 16'h213, 16'h213, 16'h2123, 16'h213, 16'h294, 16'h6aea, 16'hacd1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb1, 16'hacb0, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'ha490, 16'h8bad, 16'h3964, 16'h20c2, 16'h20c2, 16'h20c2, 16'h18a2, 16'h1061, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h83ab, 16'h8bcc, 16'h8bcc, 16'h8bcc, 16'h8bec, 16'h8bec, 16'h8bed, 16'h8cc, 16'h94c, 16'h94d, 16'h942d, 16'h942e, 16'h944e, 16'h9c4e, 16'h9c6f, 16'ha48f, 16'ha4af, 16'ha4b0, 16'h9c6e, 16'h39a4, 16'h1081, 16'h860, 16'h861, 16'h880, 16'h860, 16'h2944, 16'h39a5, 16'h2944, 16'h213, 16'h20c2, 16'h18c2, 16'h18c2, 16'h18a2, 16'h18a2, 16'h18a2, 16'h20a2, 16'h18c2, 16'h18a2, 16'h18a2, 16'h18a2, 16'h18a2, 16'h18c2, 16'h18a2, 16'h881, 16'h840, 16'h860, 16'h880, 16'h1081, 16'h292, 16'h3984, 16'h2924, 16'h2923, 16'h293, 16'h2923, 16'h2924, 16'h2924, 16'h2924, 16'h2924, 16'h294, 16'h2924, 16'h2923, 16'h2923, 16'h2923, 16'h213, 16'h213, 16'h213, 16'h294, 16'h2944, 16'h2944, 16'h213, 16'h861, 16'h020, 16'h28c1, 16'h6a84, 16'h41a6, 16'h10a6, 16'h866, 16'h865, 16'h844, 16'h842, 16'h841, 16'h840, 16'h020, 16'h840, 16'h2922, 16'h292, 16'h292, 16'h292, 16'h212, 16'h20c2, 16'h20e2, 16'h292, 16'h292, 16'h292, 16'h2922, 16'h2922, 16'h213, 16'h213, 16'h212, 16'h212, 16'h20e2, 16'h18c2, 16'h18a2, 16'h1081, 16'h1061, 16'h861, 16'h840, 16'h840, 16'h840, 16'h040, 16'h040, 16'h840, 16'h841, 16'h62a9, 16'hbd32, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'h734b, 16'h2924, 16'h213, 16'h213, 16'h213, 16'h2123, 16'h214, 16'h62ca, 16'hacd0, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacd1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hac90, 16'h8bcd, 16'h3165, 16'h20e3, 16'h20c2, 16'h20c2, 16'h18a2, 16'h1061, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h83ab, 16'h8bcc, 16'h8bec, 16'h8bec, 16'h8bec, 16'h8bec, 16'h8bed, 16'h8cd, 16'h94d, 16'h942d, 16'h942d, 16'h942e, 16'h9c4e, 16'h9c6f, 16'ha48f, 16'ha48f, 16'ha4af, 16'ha4b0, 16'h9c8f, 16'h41c5, 16'h1081, 16'h860, 16'h860, 16'h860, 16'h860, 16'h18e2, 16'h39c5, 16'h3144, 16'h213, 16'h20c3, 16'h18c2, 16'h18a2, 16'h18a2, 16'h18a2, 16'h18a2, 16'h18a2, 16'h18a3, 16'h18a2, 16'h18a2, 16'h18a2, 16'h18a2, 16'h18c2, 16'h18c3, 16'h18c3, 16'h1081, 16'h840, 16'h860, 16'h1881, 16'h3123, 16'h3984, 16'h2924, 16'h2924, 16'h293, 16'h294, 16'h294, 16'h294, 16'h2924, 16'h2924, 16'h2924, 16'h2924, 16'h2924, 16'h2923, 16'h2923, 16'h293, 16'h213, 16'h213, 16'h2923, 16'h2944, 16'h2924, 16'h213, 16'h1061, 16'h020, 16'h28e1, 16'h6a63, 16'h295, 16'h866, 16'h865, 16'h845, 16'h845, 16'h864, 16'h1063, 16'h3965, 16'h49e6, 16'h3144, 16'h3963, 16'h3984, 16'h3163, 16'h3143, 16'h3143, 16'h2922, 16'h2923, 16'h2923, 16'h293, 16'h2923, 16'h2923, 16'h2923, 16'h2923, 16'h2923, 16'h2923, 16'h2923, 16'h3123, 16'h3123, 16'h3123, 16'h2943, 16'h2923, 16'h2923, 16'h2923, 16'h213, 16'h212, 16'h20e2, 16'h18c2, 16'h18a2, 16'h18a2, 16'h6aca, 16'hbd32, 16'hc533, 16'hbd33, 16'hbd32, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd32, 16'hbd32, 16'hbd12, 16'hbd12, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'ha4b0, 16'h4a27, 16'h214, 16'h214, 16'h214, 16'h2124, 16'h214, 16'h3145, 16'h73b, 16'hacd1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb1, 16'hacd0, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacd0, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb0, 16'h8bce, 16'h3965, 16'h20e2, 16'h20c2, 16'h18c2, 16'h18a2, 16'h1061, 16'h020, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h83ab, 16'h8bcc, 16'h8bec, 16'h8bec, 16'h8bec, 16'h8bed, 16'h8cd, 16'h94d, 16'h942d, 16'h942d, 16'h942d, 16'h944e, 16'h9c4e, 16'h9c6f, 16'ha48f, 16'ha4af, 16'ha4b0, 16'hacd0, 16'ha48f, 16'h41c6, 16'h1061, 16'h860, 16'h860, 16'h860, 16'h860, 16'h860, 16'h2923, 16'h41c6, 16'h3144, 16'h213, 16'h20c2, 16'h18a2, 16'h18a2, 16'h18a1, 16'h1882, 16'h18a2, 16'h18a2, 16'h18a2, 16'h18a2, 16'h18a2, 16'h18a2, 16'h18c2, 16'h18c3, 16'h18a3, 16'h1881, 16'h18c2, 16'h20e2, 16'h20a2, 16'h3123, 16'h3964, 16'h3144, 16'h2924, 16'h2924, 16'h294, 16'h294, 16'h294, 16'h2924, 16'h2924, 16'h2924, 16'h2924, 16'h2924, 16'h2923, 16'h2923, 16'h294, 16'h3164, 16'h2923, 16'h2944, 16'h2944, 16'h3164, 16'h2944, 16'h1061, 16'h020, 16'h2081, 16'h6a86, 16'h72ea, 16'h41c9, 16'h845, 16'h845, 16'h865, 16'h864, 16'h1884, 16'h73b, 16'h9c4e, 16'h62a8, 16'h4184, 16'h4184, 16'h3984, 16'h3163, 16'h3143, 16'h3142, 16'h3143, 16'h3143, 16'h213, 16'h20e2, 16'h20e2, 16'h212, 16'h292, 16'h2923, 16'h2923, 16'h2943, 16'h3143, 16'h3143, 16'h3143, 16'h3143, 16'h3144, 16'h3143, 16'h3163, 16'h3144, 16'h3163, 16'h3163, 16'h3163, 16'h3144, 16'h3164, 16'h7b2b, 16'hbd32, 16'hc553, 16'hc553, 16'hc553, 16'hc553, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'h94e, 16'h3165, 16'h2923, 16'h2123, 16'h2924, 16'h2124, 16'h294, 16'h5a69, 16'h8bce, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hb4d1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'h93ce, 16'h3965, 16'h20e3, 16'h20c2, 16'h18c2, 16'h20c2, 16'h1061, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h83ab, 16'h8bcc, 16'h8bec, 16'h8bec, 16'h8bec, 16'h8bed, 16'h8cd, 16'h94d, 16'h94d, 16'h94d, 16'h8bed, 16'h94d, 16'h944e, 16'h9c6f, 16'h9c8f, 16'ha4af, 16'ha4b0, 16'hacd0, 16'ha4af, 16'h41e6, 16'h1081, 16'h860, 16'h860, 16'h860, 16'h860, 16'h860, 16'h1081, 16'h4a27, 16'h4a27, 16'h39a6, 16'h2924, 16'h20e3, 16'h18a2, 16'h1882, 16'h1082, 16'h1082, 16'h1881, 16'h1882, 16'h1882, 16'h18a2, 16'h18a2, 16'h18c2, 16'h18a2, 16'h18a2, 16'h10a1, 16'h18a1, 16'h2923, 16'h213, 16'h2923, 16'h3144, 16'h3144, 16'h2944, 16'h2924, 16'h2924, 16'h2924, 16'h2924, 16'h2924, 16'h2924, 16'h2924, 16'h2924, 16'h2924, 16'h2924, 16'h2924, 16'h3965, 16'h4a6, 16'h2923, 16'h3164, 16'h20e2, 16'h2923, 16'h2943, 16'h1081, 16'h020, 16'h1081, 16'h5a87, 16'h838b, 16'h6aea, 16'h2946, 16'h1085, 16'h1085, 16'h1084, 16'h3166, 16'h8bac, 16'h838b, 16'h41a5, 16'h4184, 16'h4184, 16'h4184, 16'h3984, 16'h3163, 16'h3143, 16'h3143, 16'h3143, 16'h20e2, 16'h1081, 16'h1081, 16'h18a1, 16'h18a1, 16'h18c2, 16'h20c2, 16'h20e2, 16'h20e2, 16'h293, 16'h2923, 16'h2923, 16'h2943, 16'h3143, 16'h3143, 16'h3164, 16'h3163, 16'h3163, 16'h3164, 16'h3164, 16'h3984, 16'h7b4b, 16'hbd32, 16'hc553, 16'hc553, 16'hc553, 16'hc553, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb532, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'h7b2c, 16'h2924, 16'h2924, 16'h2924, 16'h2124, 16'h2124, 16'h3145, 16'h732c, 16'h9cf, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacd1, 16'hacd1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d2, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacb1, 16'h93ee, 16'h3965, 16'h20e3, 16'h20c2, 16'h20c2, 16'h20c2, 16'h1061, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h838b, 16'h8bcc, 16'h8bec, 16'h8bec, 16'h8bec, 16'h8bed, 16'h8bed, 16'h94d, 16'h94d, 16'h8bcc, 16'h7b4b, 16'h838c, 16'h942e, 16'h9c4f, 16'h9c6f, 16'ha490, 16'ha4b0, 16'hacd0, 16'ha4af, 16'h49e6, 16'h1081, 16'h860, 16'h060, 16'h860, 16'h860, 16'h860, 16'h1081, 16'h5a48, 16'h6289, 16'h41c6, 16'h3144, 16'h3965, 16'h3145, 16'h20e4, 16'h18a3, 16'h1882, 16'h1882, 16'h1882, 16'h1882, 16'h1881, 16'h18a2, 16'h18a2, 16'h18a2, 16'h18a2, 16'h10a1, 16'h1081, 16'h18e2, 16'h18c1, 16'h1081, 16'h293, 16'h3144, 16'h2924, 16'h2924, 16'h2924, 16'h2924, 16'h2924, 16'h2924, 16'h2924, 16'h2924, 16'h2924, 16'h2924, 16'h2924, 16'h3985, 16'h5a88, 16'h5a67, 16'h2923, 16'h3164, 16'h18a2, 16'h20e2, 16'h2923, 16'h1081, 16'h020, 16'h861, 16'h2924, 16'h3164, 16'h3964, 16'h3144, 16'h2924, 16'h2924, 16'h2924, 16'h3164, 16'h41c5, 16'h41c5, 16'h2923, 16'h41c4, 16'h3983, 16'h4183, 16'h4184, 16'h3963, 16'h2922, 16'h3143, 16'h3143, 16'h20c2, 16'h1041, 16'h1061, 16'h1061, 16'h1081, 16'h1081, 16'h1081, 16'h1081, 16'h1081, 16'h1081, 16'h18a1, 16'h18a1, 16'h18c1, 16'h20c2, 16'h20e2, 16'h293, 16'h2923, 16'h2923, 16'h3143, 16'h3163, 16'h3984, 16'h7b4b, 16'hbd32, 16'hc553, 16'hc553, 16'hc553, 16'hc553, 16'hc553, 16'hc553, 16'hc553, 16'hc553, 16'hc553, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hb512, 16'hb532, 16'hb532, 16'hb512, 16'hb512, 16'hb512, 16'hb4f1, 16'h628a, 16'h2924, 16'h2924, 16'h2924, 16'h2124, 16'h2924, 16'h41a7, 16'h628a, 16'h9c4f, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d2, 16'hb4d2, 16'hb4d1, 16'hacd1, 16'hacb1, 16'h93ee, 16'h3985, 16'h20e2, 16'h20c2, 16'h20c2, 16'h20c2, 16'h1081, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h83ab, 16'h83cb, 16'h8bec, 16'h8bec, 16'h8bec, 16'h8bed, 16'h8bed, 16'h8cd, 16'h94d, 16'h83ac, 16'h732a, 16'h7b6b, 16'h94e, 16'h9c4e, 16'h942e, 16'h9c6f, 16'ha48f, 16'ha4b0, 16'ha4af, 16'h4a6, 16'h1081, 16'h860, 16'h860, 16'h860, 16'h860, 16'h860, 16'h1081, 16'h5a68, 16'h5a68, 16'h3984, 16'h1061, 16'h18a2, 16'h213, 16'h2944, 16'h3165, 16'h3144, 16'h294, 16'h20e3, 16'h18a2, 16'h18a2, 16'h18a2, 16'h10a2, 16'h10a2, 16'h10a2, 16'h1081, 16'h861, 16'h881, 16'h860, 16'h860, 16'h213, 16'h3164, 16'h2944, 16'h2924, 16'h3985, 16'h41c6, 16'h294, 16'h3165, 16'h3985, 16'h3985, 16'h3965, 16'h3144, 16'h3124, 16'h5248, 16'h73a, 16'h5247, 16'h3144, 16'h3164, 16'h18a2, 16'h1081, 16'h212, 16'h1081, 16'h020, 16'h840, 16'h293, 16'h2923, 16'h2923, 16'h3124, 16'h3124, 16'h3124, 16'h3124, 16'h2924, 16'h20e2, 16'h3144, 16'h292, 16'h39a4, 16'h3983, 16'h3983, 16'h3983, 16'h3983, 16'h3963, 16'h3963, 16'h3984, 16'h3143, 16'h2923, 16'h2922, 16'h293, 16'h292, 16'h292, 16'h20e2, 16'h20c2, 16'h1081, 16'h1061, 16'h1061, 16'h1061, 16'h1061, 16'h1061, 16'h1061, 16'h1081, 16'h18a1, 16'h18a1, 16'h18c2, 16'h20e2, 16'h2923, 16'h73b, 16'hbd33, 16'hc553, 16'hc553, 16'hc553, 16'hc553, 16'hc553, 16'hc553, 16'hc553, 16'hc553, 16'hc553, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hb532, 16'hbd32, 16'hbd32, 16'hb512, 16'hb512, 16'hacb1, 16'h5228, 16'h2924, 16'h2924, 16'h2924, 16'h2124, 16'h2924, 16'h4227, 16'h5a89, 16'hacb1, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d2, 16'hb4f2, 16'hb4f1, 16'hb4d1, 16'hacd1, 16'h93ee, 16'h3985, 16'h20e2, 16'h20c2, 16'h20c2, 16'h20c1, 16'h1081, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h7b8b, 16'h83ab, 16'h8bcc, 16'h8bec, 16'h8bec, 16'h8bec, 16'h8bec, 16'h8cc, 16'h94d, 16'h8bcc, 16'h7b6b, 16'h838c, 16'h94d, 16'h942e, 16'h942e, 16'h9c4f, 16'ha48f, 16'ha4b0, 16'ha4af, 16'h4a6, 16'h1081, 16'h860, 16'h860, 16'h860, 16'h860, 16'h860, 16'h1082, 16'h5a48, 16'h5248, 16'h3164, 16'h861, 16'h861, 16'h840, 16'h860, 16'h18a1, 16'h20e3, 16'h2923, 16'h3164, 16'h3144, 16'h2944, 16'h213, 16'h20e3, 16'h18c2, 16'h18a2, 16'h1081, 16'h861, 16'h860, 16'h860, 16'h860, 16'h2123, 16'h39a5, 16'h3165, 16'h5a69, 16'h8bad, 16'h7b4b, 16'h49e7, 16'h5a48, 16'h6268, 16'h5a68, 16'h5227, 16'h49c6, 16'h41a5, 16'h6aa9, 16'h73a, 16'h49e6, 16'h3984, 16'h3164, 16'h18a2, 16'h18a2, 16'h20e3, 16'h1081, 16'h020, 16'h840, 16'h20e2, 16'h293, 16'h293, 16'h293, 16'h2923, 16'h2923, 16'h2924, 16'h2924, 16'h2924, 16'h41c5, 16'h293, 16'h39a4, 16'h3983, 16'h3984, 16'h3983, 16'h41a4, 16'h41c4, 16'h41c4, 16'h41a4, 16'h2943, 16'h20e2, 16'h18c1, 16'h18a1, 16'h18a1, 16'h18c1, 16'h20e1, 16'h2923, 16'h2943, 16'h2923, 16'h18c2, 16'h1081, 16'h1081, 16'h1081, 16'h1081, 16'h1081, 16'h1081, 16'h1081, 16'h18a1, 16'h18a1, 16'h18c2, 16'h72ea, 16'hc553, 16'hc553, 16'hc553, 16'hc553, 16'hc553, 16'hc553, 16'hc553, 16'hc553, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hb512, 16'hacb1, 16'h4a7, 16'h2124, 16'h2924, 16'h2124, 16'h2124, 16'h3164, 16'h41e6, 16'h732b, 16'hb4f1, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4f1, 16'hb4f1, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4d2, 16'hb4d1, 16'h94e, 16'h3985, 16'h20e2, 16'h20e2, 16'h20c2, 16'h20c2, 16'h1081, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h7b6a, 16'h83ab, 16'h8bcc, 16'h8bcc, 16'h8bcc, 16'h8bcc, 16'h8bec, 16'h8cc, 16'h94d, 16'h942d, 16'h942e, 16'h942e, 16'h942e, 16'h942e, 16'h9c4f, 16'h9c6f, 16'ha48f, 16'ha4b0, 16'ha48f, 16'h4a6, 16'h1081, 16'h860, 16'h860, 16'h860, 16'h860, 16'h860, 16'h10a1, 16'h5a68, 16'h5247, 16'h3164, 16'h860, 16'h860, 16'h040, 16'h040, 16'h860, 16'h860, 16'h860, 16'h881, 16'h10a1, 16'h20e2, 16'h2923, 16'h2923, 16'h2924, 16'h293, 16'h18c2, 16'h1081, 16'h860, 16'h860, 16'h860, 16'h2924, 16'h4a8, 16'h6aca, 16'h9c50, 16'hacb0, 16'h8bad, 16'h834c, 16'h7ba, 16'h6289, 16'h5a48, 16'h527, 16'h49c6, 16'h4185, 16'h5a68, 16'h6ae9, 16'h4a7, 16'h49e6, 16'h3164, 16'h20e2, 16'h20e2, 16'h293, 16'h1081, 16'h020, 16'h841, 16'h2923, 16'h3164, 16'h3164, 16'h3164, 16'h3984, 16'h3984, 16'h3985, 16'h3165, 16'h41c6, 16'h5247, 16'h2923, 16'h39a4, 16'h3983, 16'h41a4, 16'h41c4, 16'h41a4, 16'h3984, 16'h3163, 16'h3963, 16'h212, 16'h1881, 16'h1081, 16'h1081, 16'h1081, 16'h1081, 16'h1081, 16'h1081, 16'h18a1, 16'h293, 16'h3164, 16'h2923, 16'h18a1, 16'h18a2, 16'h18a2, 16'h18a2, 16'h18c1, 16'h18c2, 16'h18c2, 16'h20c2, 16'h20e2, 16'h73a, 16'hc553, 16'hc553, 16'hc553, 16'hc553, 16'hc553, 16'hc573, 16'hc573, 16'hc573, 16'hc553, 16'hc553, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hacb1, 16'h4a8, 16'h2124, 16'h2124, 16'h2123, 16'h2124, 16'h3185, 16'h4a7, 16'h9c4f, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hb4d1, 16'hacd1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4f1, 16'hb4f1, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f2, 16'hb4d2, 16'h942f, 16'h3985, 16'h20e2, 16'h20e2, 16'h20c2, 16'h18c2, 16'h1081, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h7b6a, 16'h838b, 16'h83ab, 16'h83ab, 16'h83cb, 16'h83cc, 16'h83ec, 16'h8bec, 16'h8bed, 16'h942d, 16'h942e, 16'h94e, 16'h942e, 16'h9c4e, 16'h9c6f, 16'h9c6f, 16'h9c8f, 16'ha4af, 16'h9c8f, 16'h4a6, 16'h1081, 16'h860, 16'h860, 16'h860, 16'h860, 16'h860, 16'h18a1, 16'h5a68, 16'h4a7, 16'h2944, 16'h860, 16'h860, 16'h040, 16'h860, 16'h860, 16'h860, 16'h860, 16'h860, 16'h860, 16'h840, 16'h840, 16'h860, 16'h1061, 16'h1081, 16'h1081, 16'h840, 16'h840, 16'h860, 16'h860, 16'h2924, 16'h62aa, 16'h94f, 16'hacd1, 16'ha490, 16'h836c, 16'h834c, 16'h834b, 16'h72ea, 16'h62a9, 16'h527, 16'h49c6, 16'h3985, 16'h4a6, 16'h6ac9, 16'h4a7, 16'h4a6, 16'h3984, 16'h3985, 16'h3985, 16'h3164, 16'h18a2, 16'h840, 16'h861, 16'h3985, 16'h41c6, 16'h41a5, 16'h41a5, 16'h41a5, 16'h49c6, 16'h49e6, 16'h49e7, 16'h5227, 16'h49e6, 16'h292, 16'h3984, 16'h41c5, 16'h41a5, 16'h3963, 16'h3163, 16'h3163, 16'h3163, 16'h3163, 16'h2923, 16'h1881, 16'h1881, 16'h1881, 16'h1081, 16'h1081, 16'h1081, 16'h1081, 16'h1881, 16'h1881, 16'h20c2, 16'h3164, 16'h3144, 16'h1881, 16'h18a2, 16'h18a2, 16'h18a2, 16'h18c2, 16'h18c2, 16'h20e2, 16'h213, 16'h73b, 16'hc573, 16'hc574, 16'hc574, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc553, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hacd1, 16'h5229, 16'h2924, 16'h2124, 16'h2124, 16'h2944, 16'h3165, 16'h6aea, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'h9c2f, 16'h3985, 16'h20e2, 16'h20c2, 16'h20c2, 16'h20a2, 16'h1081, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h734a, 16'h7b6a, 16'h838b, 16'h83ab, 16'h83ab, 16'h83ac, 16'h83cc, 16'h83cc, 16'h8bec, 16'h8cd, 16'h8bed, 16'h8bed, 16'h8bed, 16'h94e, 16'h9c4e, 16'h9c4f, 16'h9c6e, 16'h9c8f, 16'h9c6e, 16'h4a6, 16'h1081, 16'h860, 16'h860, 16'h860, 16'h860, 16'h860, 16'h10a1, 16'h5a68, 16'h41e6, 16'h2923, 16'h860, 16'h860, 16'h060, 16'h060, 16'h860, 16'h860, 16'h860, 16'h860, 16'h860, 16'h860, 16'h860, 16'h860, 16'h840, 16'h840, 16'h840, 16'h040, 16'h840, 16'h840, 16'h840, 16'h18a2, 16'h7b4c, 16'hacd1, 16'hacb1, 16'ha470, 16'h7b4b, 16'h834c, 16'h836c, 16'h7b2b, 16'h6aa9, 16'h526, 16'h49c6, 16'h4185, 16'h4a6, 16'h6ac9, 16'h4a7, 16'h4a6, 16'h41c5, 16'h4a6, 16'h4a6, 16'h39a5, 16'h18a2, 16'h840, 16'h861, 16'h39a5, 16'h4a7, 16'h4a6, 16'h49e6, 16'h49c6, 16'h49e6, 16'h5227, 16'h5a47, 16'h5a68, 16'h3964, 16'h28e2, 16'h49e5, 16'h41c4, 16'h3143, 16'h3143, 16'h3143, 16'h3143, 16'h3143, 16'h3163, 16'h3984, 16'h20e2, 16'h1881, 16'h1881, 16'h1881, 16'h1081, 16'h1081, 16'h1881, 16'h1081, 16'h1081, 16'h1081, 16'h18a1, 16'h3984, 16'h2923, 16'h1881, 16'h1881, 16'h1881, 16'h18a1, 16'h18a2, 16'h18c2, 16'h20e3, 16'h73b, 16'hc573, 16'hcd74, 16'hcd74, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc573, 16'hc573, 16'hc573, 16'hc553, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd32, 16'hb4f2, 16'h6aeb, 16'h2945, 16'h2924, 16'h2965, 16'h3145, 16'h5228, 16'ha470, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d2, 16'hb4d1, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'h9c2f, 16'h3985, 16'h20e3, 16'h20c3, 16'h20c2, 16'h18c2, 16'h1081, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h7329, 16'h7b4a, 16'h7b8a, 16'h838b, 16'h838b, 16'h838c, 16'h83ac, 16'h83ac, 16'h83cc, 16'h8bec, 16'h8bec, 16'h8bed, 16'h8cd, 16'h94d, 16'h942e, 16'h944e, 16'h9c4e, 16'h9c6f, 16'h944e, 16'h4a6, 16'h861, 16'h060, 16'h860, 16'h860, 16'h860, 16'h860, 16'h10a1, 16'h5a68, 16'h41c6, 16'h2123, 16'h840, 16'h860, 16'h860, 16'h060, 16'h060, 16'h860, 16'h860, 16'h860, 16'h860, 16'h860, 16'h860, 16'h860, 16'h860, 16'h860, 16'h840, 16'h040, 16'h840, 16'h860, 16'h840, 16'h41a6, 16'h9c70, 16'hacd1, 16'hacb1, 16'h9c4f, 16'h7b2b, 16'h834b, 16'h836c, 16'h834b, 16'h6ac9, 16'h527, 16'h49c6, 16'h41a5, 16'h4a7, 16'h6ac9, 16'h526, 16'h49e6, 16'h41c5, 16'h49e5, 16'h41a5, 16'h3984, 16'h18c2, 16'h840, 16'h861, 16'h3985, 16'h4a6, 16'h5227, 16'h5a48, 16'h527, 16'h49e6, 16'h4a6, 16'h5227, 16'h5247, 16'h41c5, 16'h41c5, 16'h49e5, 16'h3123, 16'h2922, 16'h2922, 16'h2922, 16'h2923, 16'h3143, 16'h3143, 16'h3143, 16'h2923, 16'h1881, 16'h1881, 16'h1881, 16'h1081, 16'h1081, 16'h1081, 16'h1081, 16'h1081, 16'h1081, 16'h1081, 16'h20e3, 16'h3985, 16'h18a2, 16'h1081, 16'h1081, 16'h1881, 16'h1881, 16'h18a1, 16'h20e3, 16'h73b, 16'hc573, 16'hcd94, 16'hcd94, 16'hcd74, 16'hcd74, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc573, 16'hc573, 16'hc573, 16'hc553, 16'hc553, 16'hc553, 16'hc553, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd32, 16'h8bce, 16'h41a7, 16'h5229, 16'h41c7, 16'h41c7, 16'h8bce, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f2, 16'hb4f1, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'h9c4f, 16'h3985, 16'h20e3, 16'h20c2, 16'h20c2, 16'h20c2, 16'h1081, 16'h020, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h7329, 16'h734a, 16'h7b6a, 16'h7b6a, 16'h7b6b, 16'h7b6b, 16'h838b, 16'h83ab, 16'h83ac, 16'h83cc, 16'h83cc, 16'h8bec, 16'h8bed, 16'h8cd, 16'h942d, 16'h942e, 16'h942e, 16'h83ac, 16'h7b6a, 16'h41e5, 16'h860, 16'h060, 16'h860, 16'h860, 16'h860, 16'h860, 16'h18a1, 16'h5a68, 16'h39c6, 16'h213, 16'h840, 16'h860, 16'h060, 16'h860, 16'h860, 16'h860, 16'h860, 16'h860, 16'h860, 16'h860, 16'h860, 16'h860, 16'h860, 16'h860, 16'h040, 16'h040, 16'h840, 16'h860, 16'h1881, 16'h7b4c, 16'hb4d2, 16'hacb1, 16'ha470, 16'h9c4f, 16'h7b2b, 16'h836c, 16'h838c, 16'h834b, 16'h72c9, 16'h527, 16'h49c6, 16'h41c6, 16'h4a27, 16'h6ae9, 16'h5227, 16'h4a7, 16'h41a5, 16'h41a5, 16'h3164, 16'h3164, 16'h18c2, 16'h840, 16'h861, 16'h3985, 16'h49e6, 16'h5247, 16'h6289, 16'h5247, 16'h49e6, 16'h4a6, 16'h4a6, 16'h5227, 16'h49c6, 16'h5227, 16'h3984, 16'h292, 16'h2923, 16'h3122, 16'h3143, 16'h3143, 16'h3163, 16'h3163, 16'h292, 16'h293, 16'h18a1, 16'h1881, 16'h1081, 16'h1881, 16'h1881, 16'h1881, 16'h1081, 16'h1081, 16'h1081, 16'h1081, 16'h1081, 16'h3985, 16'h3144, 16'h1081, 16'h1061, 16'h1081, 16'h1081, 16'h1882, 16'h20c3, 16'h73b, 16'hc574, 16'hcd94, 16'hcd94, 16'hcd94, 16'hcd94, 16'hcd94, 16'hcd94, 16'hcd94, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc573, 16'hc573, 16'hc573, 16'hc553, 16'hc553, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd33, 16'hbd33, 16'hb4f2, 16'h836d, 16'h6aab, 16'h6269, 16'h8bce, 16'hbd12, 16'hbd12, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f2, 16'hb4f1, 16'hb4f2, 16'hb4f1, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'h9c50, 16'h3985, 16'h20e3, 16'h20e2, 16'h20c2, 16'h20c2, 16'h1061, 16'h020, 16'h020, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h6b9, 16'h6b29, 16'h734a, 16'h734a, 16'h7b4a, 16'h7b6b, 16'h7b6b, 16'h838b, 16'h838b, 16'h83ab, 16'h83ac, 16'h83cc, 16'h8bec, 16'h8bed, 16'h8cd, 16'h942d, 16'h8cd, 16'h5227, 16'h20c2, 16'h18c1, 16'h860, 16'h860, 16'h860, 16'h860, 16'h860, 16'h860, 16'h10a1, 16'h5248, 16'h39a6, 16'h213, 16'h860, 16'h860, 16'h860, 16'h860, 16'h860, 16'h860, 16'h860, 16'h860, 16'h860, 16'h860, 16'h860, 16'h860, 16'h860, 16'h860, 16'h040, 16'h040, 16'h840, 16'h860, 16'h3965, 16'ha470, 16'hb4f2, 16'hacb1, 16'ha470, 16'h9c2f, 16'h7b2b, 16'h836c, 16'h8b8c, 16'h834c, 16'h6aca, 16'h527, 16'h49e6, 16'h49c6, 16'h5227, 16'h6ae9, 16'h5227, 16'h4a7, 16'h41c6, 16'h4a6, 16'h41a5, 16'h3985, 16'h18a2, 16'h840, 16'h861, 16'h39a5, 16'h49e6, 16'h4a6, 16'h5227, 16'h5227, 16'h4a6, 16'h4a6, 16'h4a6, 16'h4a7, 16'h49c6, 16'h5247, 16'h41a5, 16'h3143, 16'h3163, 16'h3163, 16'h3143, 16'h3143, 16'h3163, 16'h3163, 16'h293, 16'h20e2, 16'h20c2, 16'h1081, 16'h1081, 16'h1081, 16'h1081, 16'h1081, 16'h1081, 16'h1081, 16'h1081, 16'h1081, 16'h1081, 16'h293, 16'h39a5, 16'h1081, 16'h1061, 16'h1081, 16'h1081, 16'h1081, 16'h18a2, 16'h73b, 16'hcd94, 16'hcd94, 16'hcd94, 16'hcd94, 16'hcd94, 16'hcd94, 16'hcd94, 16'hcd94, 16'hcd94, 16'hcd94, 16'hcd74, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc573, 16'hc553, 16'hc553, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd33, 16'hbd32, 16'hbd32, 16'hacb1, 16'hb4d2, 16'hbd32, 16'hbd32, 16'hbd12, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f2, 16'hb4f1, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4f1, 16'hb4d1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb512, 16'hb4f2, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'h9c50, 16'h3985, 16'h20e3, 16'h20e2, 16'h20c2, 16'h20c2, 16'h1061, 16'h020, 16'h020, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h62e8, 16'h6b9, 16'h7329, 16'h732a, 16'h7329, 16'h734a, 16'h7b4a, 16'h7b6b, 16'h7b6b, 16'h7b8b, 16'h838b, 16'h83ac, 16'h83cc, 16'h8bcc, 16'h8bed, 16'h8cd, 16'h8cd, 16'h4a26, 16'h1081, 16'h1081, 16'h860, 16'h860, 16'h840, 16'h860, 16'h860, 16'h060, 16'h1081, 16'h5268, 16'h39a5, 16'h213, 16'h860, 16'h860, 16'h060, 16'h060, 16'h060, 16'h860, 16'h860, 16'h860, 16'h860, 16'h860, 16'h860, 16'h860, 16'h860, 16'h860, 16'h040, 16'h020, 16'h840, 16'h1061, 16'h6acb, 16'hb4f2, 16'hb4d1, 16'hacd1, 16'ha470, 16'h9c2f, 16'h7bb, 16'h836c, 16'h8b8c, 16'h834c, 16'h6aa9, 16'h526, 16'h49e6, 16'h49c6, 16'h5227, 16'h6ae9, 16'h5227, 16'h49e6, 16'h41c5, 16'h5247, 16'h5227, 16'h41c6, 16'h18c2, 16'h840, 16'h841, 16'h3144, 16'h39a5, 16'h4a6, 16'h5247, 16'h5227, 16'h4a6, 16'h4a6, 16'h49e6, 16'h5227, 16'h49c6, 16'h5227, 16'h5226, 16'h3984, 16'h3963, 16'h3163, 16'h3163, 16'h3143, 16'h3143, 16'h3163, 16'h292, 16'h20e2, 16'h292, 16'h1081, 16'h1081, 16'h1081, 16'h1081, 16'h1081, 16'h1081, 16'h1081, 16'h1081, 16'h1081, 16'h1081, 16'h20c2, 16'h39a5, 16'h1081, 16'h1061, 16'h1061, 16'h1081, 16'h1081, 16'h18a2, 16'h73b, 16'hcd94, 16'hcdb5, 16'hcdb4, 16'hcdb4, 16'hcd94, 16'hcd95, 16'hcd94, 16'hcd94, 16'hcd94, 16'hcd94, 16'hcd74, 16'hcd74, 16'hcd74, 16'hc574, 16'hc574, 16'hc574, 16'hc573, 16'hc573, 16'hc553, 16'hc553, 16'hc553, 16'hc553, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hacd1, 16'hb4d1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb512, 16'hb4f2, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hbd12, 16'hbd12, 16'hb4f2, 16'ha471, 16'h3986, 16'h20e3, 16'h20e2, 16'h20c2, 16'h20c2, 16'h1061, 16'h020, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h5aa8, 16'h62c8, 16'h6ae9, 16'h6ae9, 16'h6b9, 16'h6b29, 16'h732a, 16'h734a, 16'h7b4a, 16'h7b6b, 16'h7b6b, 16'h7b8c, 16'h83ac, 16'h83cc, 16'h83cc, 16'h8bec, 16'h8bec, 16'h5246, 16'h18a1, 16'h1081, 16'h860, 16'h860, 16'h860, 16'h060, 16'h860, 16'h060, 16'h1081, 16'h5247, 16'h3185, 16'h20e3, 16'h860, 16'h860, 16'h060, 16'h060, 16'h060, 16'h060, 16'h060, 16'h060, 16'h860, 16'h860, 16'h060, 16'h860, 16'h860, 16'h860, 16'h040, 16'h040, 16'h10a2, 16'h5228, 16'ha470, 16'hb4f2, 16'hb4d1, 16'hacd1, 16'ha46f, 16'h9ce, 16'h7bb, 16'h838c, 16'h8b8c, 16'h834c, 16'h6aa9, 16'h5226, 16'h4a6, 16'h49e6, 16'h527, 16'h6aea, 16'h5227, 16'h49c6, 16'h41a5, 16'h5247, 16'h5a68, 16'h5228, 16'h20c3, 16'h840, 16'h841, 16'h3164, 16'h3143, 16'h3984, 16'h41a5, 16'h41c5, 16'h41c5, 16'h49c5, 16'h49e5, 16'h4a6, 16'h41c5, 16'h4a6, 16'h5226, 16'h3984, 16'h3964, 16'h3963, 16'h3163, 16'h3163, 16'h3964, 16'h3163, 16'h20c2, 16'h18c1, 16'h2923, 16'h1060, 16'h860, 16'h860, 16'h860, 16'h1060, 16'h1060, 16'h1061, 16'h1061, 16'h1081, 16'h1081, 16'h20c2, 16'h3984, 16'h1061, 16'h1061, 16'h1061, 16'h1081, 16'h1081, 16'h18a2, 16'h73b, 16'hcdb4, 16'hd5b5, 16'hcdb5, 16'hcdb5, 16'hcdb5, 16'hcd95, 16'hcd95, 16'hcd95, 16'hcd94, 16'hcd94, 16'hcd94, 16'hcd94, 16'hcd74, 16'hcd74, 16'hcd74, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc573, 16'hc554, 16'hc553, 16'hc553, 16'hc553, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hb512, 16'ha491, 16'h3986, 16'h20e2, 16'h20e2, 16'h20c2, 16'h20c2, 16'h1081, 16'h020, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h5a87, 16'h5a88, 16'h62a8, 16'h62c8, 16'h6ac9, 16'h6ae9, 16'h6ae9, 16'h6b9, 16'h732a, 16'h734a, 16'h736a, 16'h7b6b, 16'h7b8b, 16'h83ab, 16'h83cc, 16'h83cc, 16'h8bcc, 16'h5246, 16'h10a1, 16'h860, 16'h860, 16'h860, 16'h860, 16'h860, 16'h860, 16'h860, 16'h1081, 16'h4a27, 16'h3164, 16'h18c2, 16'h840, 16'h860, 16'h040, 16'h060, 16'h060, 16'h060, 16'h860, 16'h840, 16'h840, 16'h860, 16'h860, 16'h860, 16'h860, 16'h860, 16'h040, 16'h840, 16'h20e3, 16'h8bad, 16'hbd32, 16'hb4f2, 16'hb4d1, 16'hacb0, 16'ha46f, 16'h9c2e, 16'h7bb, 16'h8b8c, 16'h8bac, 16'h836c, 16'h6ac9, 16'h5227, 16'h4a7, 16'h49e6, 16'h4a6, 16'h6aea, 16'h5227, 16'h4a6, 16'h49e6, 16'h5247, 16'h5227, 16'h5248, 16'h20e3, 16'h840, 16'h1081, 16'h4a26, 16'h4a6, 16'h3164, 16'h3964, 16'h3984, 16'h41a5, 16'h41c5, 16'h49e5, 16'h4a6, 16'h41a5, 16'h3964, 16'h49e5, 16'h4184, 16'h3964, 16'h3963, 16'h3163, 16'h3163, 16'h3163, 16'h3963, 16'h20c2, 16'h1061, 16'h2923, 16'h1081, 16'h840, 16'h840, 16'h860, 16'h860, 16'h860, 16'h840, 16'h860, 16'h1060, 16'h1060, 16'h2923, 16'h2943, 16'h1060, 16'h1060, 16'h1060, 16'h1061, 16'h1081, 16'h18a2, 16'h73b, 16'hcdb4, 16'hd5b5, 16'hd5b5, 16'hd5b5, 16'hcdb5, 16'hcdb5, 16'hcdb5, 16'hcdb5, 16'hcdb4, 16'hcd94, 16'hcd94, 16'hcd94, 16'hcd94, 16'hcd94, 16'hcd74, 16'hcd74, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc573, 16'hc573, 16'hc573, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'ha491, 16'h3986, 16'h20e3, 16'h20e2, 16'h20c2, 16'h20c2, 16'h1081, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h62a7, 16'h62a8, 16'h62c8, 16'h62c8, 16'h62c8, 16'h6ae8, 16'h6ae8, 16'h6b9, 16'h6b9, 16'h6b9, 16'h7329, 16'h734a, 16'h736a, 16'h7b6b, 16'h7b8b, 16'h83ab, 16'h83ac, 16'h4a46, 16'h10a1, 16'h860, 16'h860, 16'h860, 16'h860, 16'h060, 16'h060, 16'h060, 16'h1081, 16'h4a27, 16'h2944, 16'h10a2, 16'h840, 16'h840, 16'h040, 16'h040, 16'h060, 16'h040, 16'h060, 16'h060, 16'h860, 16'h860, 16'h860, 16'h860, 16'h860, 16'h860, 16'h840, 16'h840, 16'h294, 16'h9c70, 16'hbd53, 16'hb512, 16'hb4d1, 16'hacb0, 16'ha470, 16'h94e, 16'h72ea, 16'h8bad, 16'h8bac, 16'h836c, 16'h6ac9, 16'h5227, 16'h4a7, 16'h49e6, 16'h4a7, 16'h6aea, 16'h527, 16'h4a6, 16'h4a6, 16'h5248, 16'h4a6, 16'h5247, 16'h20e3, 16'h840, 16'h840, 16'h3985, 16'h5a88, 16'h5227, 16'h41c5, 16'h41c5, 16'h41c5, 16'h41c5, 16'h49e6, 16'h4a6, 16'h41c5, 16'h3964, 16'h49e5, 16'h3984, 16'h3984, 16'h3983, 16'h3963, 16'h3143, 16'h3143, 16'h3163, 16'h20e2, 16'h1061, 16'h2923, 16'h18a1, 16'h840, 16'h840, 16'h840, 16'h840, 16'h840, 16'h840, 16'h840, 16'h860, 16'h1081, 16'h3164, 16'h18a1, 16'h860, 16'h860, 16'h860, 16'h1060, 16'h1061, 16'h18a2, 16'h73b, 16'hcdb5, 16'hd5d5, 16'hd5d5, 16'hd5b5, 16'hd5b5, 16'hd5b5, 16'hcdb5, 16'hcdb5, 16'hcdb5, 16'hcdb4, 16'hcdb4, 16'hcd94, 16'hcd94, 16'hcd94, 16'hcd94, 16'hcd94, 16'hcd94, 16'hcd94, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc573, 16'hc573, 16'hc573, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd52, 16'hbd32, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f2, 16'hb4f1, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hbd12, 16'hb512, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd32, 16'hbd12, 16'hbd12, 16'ha491, 16'h3986, 16'h20e3, 16'h20c2, 16'h20c2, 16'h18c2, 16'h1061, 16'h020, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h62c8, 16'h62c8, 16'h62c9, 16'h6ae9, 16'h6ae9, 16'h6ae9, 16'h6b9, 16'h6b29, 16'h6b29, 16'h7329, 16'h734a, 16'h734a, 16'h736a, 16'h7b6b, 16'h7b8b, 16'h838b, 16'h838b, 16'h4a46, 16'h10c1, 16'h860, 16'h860, 16'h860, 16'h860, 16'h860, 16'h060, 16'h860, 16'h20e2, 16'h4a27, 16'h2944, 16'h1081, 16'h840, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h860, 16'h840, 16'h860, 16'h860, 16'h860, 16'h860, 16'h840, 16'h841, 16'h41c7, 16'hb512, 16'hbd33, 16'hb4f2, 16'hacd1, 16'hacb0, 16'ha450, 16'h94e, 16'h72ca, 16'h8b8d, 16'h8bac, 16'h836c, 16'h6ac9, 16'h5227, 16'h527, 16'h49e6, 16'h5227, 16'h6aea, 16'h527, 16'h527, 16'h527, 16'h62ca, 16'h5228, 16'h5247, 16'h213, 16'h840, 16'h840, 16'h2944, 16'h41e5, 16'h5a88, 16'h5227, 16'h49e6, 16'h49e6, 16'h49e6, 16'h49e6, 16'h4a7, 16'h49e6, 16'h41c5, 16'h49e5, 16'h3984, 16'h3984, 16'h3983, 16'h3163, 16'h3143, 16'h3143, 16'h3163, 16'h20e2, 16'h1081, 16'h212, 16'h18a1, 16'h10a1, 16'h860, 16'h860, 16'h860, 16'h860, 16'h860, 16'h860, 16'h860, 16'h2943, 16'h2943, 16'h860, 16'h860, 16'h860, 16'h861, 16'h1060, 16'h1061, 16'h1881, 16'h73b, 16'hd5d5, 16'hd5d5, 16'hd5d5, 16'hd5d5, 16'hd5d5, 16'hd5d5, 16'hd5b5, 16'hd5b5, 16'hcdb5, 16'hcdb5, 16'hcdb5, 16'hcdb5, 16'hcdb4, 16'hcd94, 16'hcd94, 16'hcd94, 16'hcd94, 16'hcd94, 16'hcd74, 16'hcd74, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc573, 16'hc573, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb512, 16'hb512, 16'hbd12, 16'hb512, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hbd12, 16'ha490, 16'h3985, 16'h20e2, 16'h20e2, 16'h20c2, 16'h18c2, 16'h1081, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h62c8, 16'h62e9, 16'h6ae9, 16'h6ae9, 16'h6b9, 16'h6b9, 16'h732a, 16'h7329, 16'h7349, 16'h734a, 16'h736a, 16'h7b6b, 16'h7b8b, 16'h83ab, 16'h83ac, 16'h83ac, 16'h83cc, 16'h5266, 16'h10c1, 16'h860, 16'h860, 16'h860, 16'h860, 16'h860, 16'h060, 16'h881, 16'h2923, 16'h5247, 16'h2924, 16'h861, 16'h860, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h840, 16'h860, 16'h860, 16'h860, 16'h860, 16'h1062, 16'h73c, 16'hc553, 16'hbd32, 16'hb4f2, 16'hacd1, 16'hac90, 16'h9c4f, 16'h94e, 16'h72ea, 16'h8bad, 16'h8b8d, 16'h834c, 16'h6aa9, 16'h5227, 16'h5227, 16'h49e6, 16'h5227, 16'h72ea, 16'h527, 16'h4a7, 16'h527, 16'h6aca, 16'h62aa, 16'h5a68, 16'h213, 16'h840, 16'h840, 16'h2944, 16'h3184, 16'h5a68, 16'h6ac9, 16'h5227, 16'h5227, 16'h527, 16'h4a6, 16'h4a7, 16'h49c6, 16'h41a5, 16'h49e5, 16'h4184, 16'h3984, 16'h3963, 16'h3163, 16'h3163, 16'h3163, 16'h3163, 16'h292, 16'h20e2, 16'h292, 16'h18a1, 16'h18e2, 16'h1081, 16'h1060, 16'h860, 16'h860, 16'h860, 16'h1060, 16'h293, 16'h2943, 16'h1060, 16'h1060, 16'h860, 16'h860, 16'h1061, 16'h1061, 16'h1061, 16'h1882, 16'h73b, 16'hd5d5, 16'hd5f6, 16'hd5d5, 16'hd5d5, 16'hd5d5, 16'hd5d5, 16'hd5d5, 16'hd5d5, 16'hd5b5, 16'hd5b5, 16'hcdb5, 16'hcdb5, 16'hcdb5, 16'hcdb5, 16'hcdb4, 16'hcd94, 16'hcd94, 16'hcd94, 16'hcd94, 16'hcd74, 16'hcd74, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc573, 16'hc573, 16'hc553, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hbd12, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb512, 16'hb512, 16'hb4f2, 16'hb512, 16'hb512, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hbd12, 16'ha450, 16'h3985, 16'h20e2, 16'h20e2, 16'h20c2, 16'h18c2, 16'h1081, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h6ae9, 16'h6ae9, 16'h6b9, 16'h6b9, 16'h6b29, 16'h732a, 16'h732a, 16'h734a, 16'h736b, 16'h7b6b, 16'h7b8b, 16'h7b8b, 16'h83ac, 16'h83cc, 16'h83cc, 16'h8bcc, 16'h8bec, 16'h5287, 16'h18c1, 16'h860, 16'h860, 16'h060, 16'h060, 16'h060, 16'h060, 16'h060, 16'h881, 16'h426, 16'h18e2, 16'h840, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h840, 16'h040, 16'h840, 16'h861, 16'h20e4, 16'h9c50, 16'hc574, 16'hbd32, 16'hb4f2, 16'hb4d1, 16'hacb0, 16'h9c2f, 16'h93ee, 16'h72eb, 16'h8bcd, 16'h8b8c, 16'h834b, 16'h6aa9, 16'h5a27, 16'h5227, 16'h49e6, 16'h5227, 16'h73a, 16'h5227, 16'h4a7, 16'h4a7, 16'h62ca, 16'h73a, 16'h5a88, 16'h2923, 16'h840, 16'h840, 16'h3164, 16'h4a6, 16'h5227, 16'h6ac9, 16'h72e9, 16'h6aa9, 16'h5a47, 16'h5227, 16'h527, 16'h49e5, 16'h41a5, 16'h49e5, 16'h4184, 16'h3984, 16'h3964, 16'h3163, 16'h3163, 16'h3163, 16'h3163, 16'h20e2, 16'h20e3, 16'h18c2, 16'h18a1, 16'h20e2, 16'h20e2, 16'h18c2, 16'h18c2, 16'h18a2, 16'h18a2, 16'h2923, 16'h3144, 16'h18a1, 16'h1060, 16'h1060, 16'h1060, 16'h1060, 16'h1061, 16'h1061, 16'h1061, 16'h18a2, 16'h732b, 16'hd5f5, 16'hd5f6, 16'hd5f6, 16'hd5f6, 16'hd5f6, 16'hd5d5, 16'hd5d5, 16'hd5d5, 16'hd5d5, 16'hd5d5, 16'hd5d5, 16'hcdb5, 16'hcdb5, 16'hcdb5, 16'hcdb4, 16'hcdb5, 16'hcdb5, 16'hcd94, 16'hcd94, 16'hcd94, 16'hcd94, 16'hcd94, 16'hcd74, 16'hc574, 16'hc574, 16'hc574, 16'hc573, 16'hc573, 16'hc553, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd33, 16'hbd12, 16'hbd33, 16'hbd32, 16'ha470, 16'h3985, 16'h20e2, 16'h20e2, 16'h20c2, 16'h18c2, 16'h1081, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h6b9, 16'h6b9, 16'h6b9, 16'h732a, 16'h734a, 16'h734a, 16'h7b6b, 16'h7b6b, 16'h7b8b, 16'h7bab, 16'h83ac, 16'h83cc, 16'h83cc, 16'h8bed, 16'h8bed, 16'h8cd, 16'h8cd, 16'h5aa8, 16'h18c1, 16'h860, 16'h860, 16'h060, 16'h060, 16'h860, 16'h840, 16'h840, 16'h2123, 16'h39c5, 16'h1081, 16'h860, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h840, 16'h840, 16'h840, 16'h841, 16'h861, 16'h5229, 16'hbd33, 16'hc553, 16'hbd12, 16'hb4f2, 16'hb4d1, 16'hacb0, 16'h9c2f, 16'h93ee, 16'h73b, 16'h93cd, 16'h8b8d, 16'h834b, 16'h6aa9, 16'h5a27, 16'h5227, 16'h49e6, 16'h5227, 16'h73a, 16'h5227, 16'h4a7, 16'h49e6, 16'h6289, 16'h6288, 16'h5a68, 16'h2924, 16'h840, 16'h841, 16'h41a5, 16'h5a68, 16'h5a68, 16'h5a47, 16'h5a46, 16'h739, 16'h7b4b, 16'h6ae9, 16'h5a68, 16'h4a6, 16'h41a5, 16'h49e6, 16'h4184, 16'h3984, 16'h3963, 16'h3963, 16'h3963, 16'h3963, 16'h3963, 16'h292, 16'h20c2, 16'h840, 16'h820, 16'h841, 16'h18c2, 16'h1061, 16'h1081, 16'h212, 16'h2943, 16'h2943, 16'h2923, 16'h2923, 16'h2923, 16'h2923, 16'h20e3, 16'h18c2, 16'h1081, 16'h861, 16'h861, 16'h1882, 16'h73b, 16'hd5f6, 16'hddf6, 16'hd5f6, 16'hd5f6, 16'hd5f6, 16'hd5f6, 16'hd5f5, 16'hd5d5, 16'hd5d5, 16'hd5d5, 16'hd5d5, 16'hcdd5, 16'hcdb5, 16'hcdb5, 16'hcdb5, 16'hcdb5, 16'hcdb5, 16'hcdb5, 16'hcdb4, 16'hcd94, 16'hcd94, 16'hcd94, 16'hcd94, 16'hcd74, 16'hc574, 16'hc574, 16'hc574, 16'hc573, 16'hc573, 16'hc553, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hbd12, 16'hb512, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb512, 16'hb512, 16'hb512, 16'hbd12, 16'hb512, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd32, 16'hbd32, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd13, 16'hbd32, 16'ha490, 16'h3965, 16'h20e2, 16'h20e2, 16'h20c2, 16'h18c2, 16'h1061, 16'h020, 16'h00, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h6b9, 16'h6b29, 16'h732a, 16'h734a, 16'h736a, 16'h7b6b, 16'h7b8b, 16'h83ab, 16'h83ac, 16'h83cc, 16'h83ec, 16'h8bed, 16'h8cd, 16'h8cd, 16'h94d, 16'h942d, 16'h942d, 16'h5aa8, 16'h18c1, 16'h860, 16'h860, 16'h860, 16'h860, 16'h840, 16'h840, 16'h1082, 16'h62c9, 16'h427, 16'h1924, 16'h1081, 16'h860, 16'h860, 16'h041, 16'h860, 16'h861, 16'h840, 16'h840, 16'h840, 16'h040, 16'h040, 16'h840, 16'h840, 16'h840, 16'h841, 16'h1082, 16'h7b4d, 16'hc574, 16'hc553, 16'hb512, 16'hb4f2, 16'hacd1, 16'hacb0, 16'h9c2f, 16'h93ee, 16'h7bb, 16'h93cd, 16'h836c, 16'h7b2b, 16'h6a89, 16'h5a28, 16'h5a28, 16'h526, 16'h5227, 16'h73a, 16'h5227, 16'h527, 16'h4a6, 16'h5a48, 16'h41c5, 16'h41c5, 16'h2924, 16'h841, 16'h840, 16'h39a5, 16'h5a47, 16'h5a47, 16'h6267, 16'h6246, 16'h72e9, 16'h8bab, 16'h72c9, 16'h6aa9, 16'h5a67, 16'h5226, 16'h4a6, 16'h4184, 16'h3984, 16'h3984, 16'h3963, 16'h3963, 16'h3963, 16'h3963, 16'h3143, 16'h18a1, 16'h820, 16'h820, 16'h820, 16'h18c2, 16'h18c2, 16'h18c2, 16'h20e2, 16'h1081, 16'h860, 16'h18c1, 16'h1881, 16'h1061, 16'h18c2, 16'h293, 16'h2923, 16'h2924, 16'h293, 16'h20e3, 16'h20c3, 16'h73b, 16'hd5f6, 16'hde16, 16'hde16, 16'hd616, 16'hd616, 16'hd5f6, 16'hd5f6, 16'hd5f6, 16'hd5d5, 16'hd5d5, 16'hd5d5, 16'hd5d5, 16'hd5d5, 16'hd5d5, 16'hd5b5, 16'hcdb5, 16'hcdb5, 16'hcdb5, 16'hcdb5, 16'hcd94, 16'hcd94, 16'hcd94, 16'hcd94, 16'hc594, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc573, 16'hc573, 16'hc553, 16'hc553, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hbd12, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb512, 16'hb512, 16'hb4f2, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hbd12, 16'hbd12, 16'hb512, 16'hb512, 16'hbd12, 16'hbd12, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd33, 16'hbd32, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd33, 16'ha490, 16'h3966, 16'h20e3, 16'h20e2, 16'h20e2, 16'h20c2, 16'h1061, 16'h020, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h7329, 16'h734a, 16'h734a, 16'h7b6a, 16'h7b8b, 16'h838c, 16'h83ac, 16'h83cc, 16'h8bec, 16'h8cc, 16'h8cd, 16'h94d, 16'h942d, 16'h942d, 16'h944e, 16'h944e, 16'h942d, 16'h62e8, 16'h18c1, 16'h860, 16'h860, 16'h860, 16'h860, 16'h840, 16'h840, 16'h10a2, 16'h6b4b, 16'h4248, 16'h3228, 16'h18e3, 16'h881, 16'h882, 16'h882, 16'h2124, 16'h4a7, 16'h41c6, 16'h3985, 16'h3164, 16'h2923, 16'h861, 16'h18a2, 16'h1082, 16'h861, 16'h861, 16'h18a3, 16'h9430, 16'hc574, 16'hc554, 16'hb512, 16'hb4d2, 16'hacd1, 16'hac90, 16'h9c2f, 16'h93ee, 16'h7b2b, 16'h93cd, 16'h836c, 16'h73b, 16'h6a89, 16'h5a48, 16'h5a48, 16'h526, 16'h527, 16'h73a, 16'h5227, 16'h527, 16'h49e6, 16'h5a48, 16'h3964, 16'h3964, 16'h3164, 16'h841, 16'h840, 16'h3164, 16'h5227, 16'h5a47, 16'h5a47, 16'h526, 16'h6267, 16'h6ac9, 16'h72e9, 16'h6ac9, 16'h62a8, 16'h6ae9, 16'h6ae9, 16'h5a87, 16'h5a47, 16'h5226, 16'h526, 16'h49e5, 16'h49e5, 16'h49c5, 16'h3984, 16'h293, 16'h20e2, 16'h20e2, 16'h20e2, 16'h20e3, 16'h213, 16'h1081, 16'h840, 16'h820, 16'h840, 16'h1081, 16'h841, 16'h840, 16'h841, 16'h1061, 16'h861, 16'h861, 16'h1081, 16'h18c2, 16'h294, 16'h834c, 16'hde16, 16'hde16, 16'hde16, 16'hd616, 16'hd616, 16'hd5f6, 16'hd5f6, 16'hd5f6, 16'hd5f6, 16'hd5f5, 16'hd5f5, 16'hd5d5, 16'hd5d5, 16'hd5d5, 16'hd5d5, 16'hd5b5, 16'hcdb5, 16'hcdb5, 16'hcdb5, 16'hcdb5, 16'hcd94, 16'hcd94, 16'hcd94, 16'hcd94, 16'hc594, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc573, 16'hc573, 16'hc573, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hbd12, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hbd12, 16'hbd12, 16'hbd32, 16'hbd12, 16'hbd13, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd33, 16'ha470, 16'h3965, 16'h20e3, 16'h20e2, 16'h20c2, 16'h20c2, 16'h1061, 16'h020, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h734a, 16'h736a, 16'h7b8b, 16'h7b8b, 16'h83ab, 16'h83cc, 16'h8bec, 16'h8cd, 16'h8cd, 16'h942d, 16'h942d, 16'h944e, 16'h944e, 16'h944e, 16'h944e, 16'h946e, 16'h944e, 16'h6ae9, 16'h18c1, 16'h860, 16'h860, 16'h060, 16'h860, 16'h860, 16'h860, 16'h10a2, 16'h6b4b, 16'h4248, 16'h3a27, 16'h193, 16'h8a1, 16'h8a2, 16'h8a2, 16'h2964, 16'h739, 16'h7b2a, 16'h7b2a, 16'h836a, 16'h732a, 16'h20e3, 16'h5a68, 16'h5a89, 16'h2966, 16'h2125, 16'h3967, 16'hacb2, 16'hc574, 16'hc554, 16'hbd32, 16'hb4d1, 16'hacb1, 16'ha490, 16'h9c4f, 16'h93ed, 16'h7b2b, 16'h93ce, 16'h8b8c, 16'h7ba, 16'h6aa9, 16'h6268, 16'h5a48, 16'h49e7, 16'h527, 16'h73a, 16'h5227, 16'h527, 16'h49e6, 16'h5a67, 16'h3964, 16'h3984, 16'h3185, 16'h841, 16'h020, 16'h18c2, 16'h3143, 16'h49c4, 16'h5226, 16'h3984, 16'h49e5, 16'h5226, 16'h6aa9, 16'h6289, 16'h527, 16'h49c6, 16'h4a6, 16'h41a4, 16'h4184, 16'h4184, 16'h3984, 16'h3984, 16'h3984, 16'h3984, 16'h3143, 16'h292, 16'h212, 16'h20e2, 16'h20c2, 16'h18a1, 16'h20e3, 16'h18a2, 16'h1081, 16'h1081, 16'h18a1, 16'h18c2, 16'h18a2, 16'h18a2, 16'h18c2, 16'h18c2, 16'h20e2, 16'h20e2, 16'h18c2, 16'h20c2, 16'h20e3, 16'h7b4c, 16'hde16, 16'hde16, 16'hde16, 16'hde16, 16'hde16, 16'hd616, 16'hd616, 16'hd5f6, 16'hd5f6, 16'hd5f6, 16'hd5f5, 16'hd5f5, 16'hd5d5, 16'hd5d5, 16'hd5d5, 16'hd5d5, 16'hd5d5, 16'hcdb5, 16'hcdb5, 16'hcdb5, 16'hcdb5, 16'hcdb4, 16'hcd94, 16'hcd94, 16'hcd94, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc553, 16'hc553, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hbd12, 16'hbd12, 16'hbd32, 16'hbd12, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd33, 16'ha470, 16'h3965, 16'h20e2, 16'h20e2, 16'h20c2, 16'h20c2, 16'h1081, 16'h020, 16'h020, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h736a, 16'h7b8b, 16'h83ac, 16'h83cc, 16'h8bec, 16'h8cd, 16'h8cd, 16'h942d, 16'h942e, 16'h944e, 16'h944e, 16'h9c4f, 16'h9c6f, 16'h9c6e, 16'h9c6f, 16'h9c6e, 16'h9c6e, 16'h6b9, 16'h18e1, 16'h860, 16'h840, 16'h881, 16'h2944, 16'h18c2, 16'h10a1, 16'h10a2, 16'h4a67, 16'h31e6, 16'h31e6, 16'h193, 16'h881, 16'h8a2, 16'h8a2, 16'h3164, 16'h739, 16'h7b4a, 16'h7b4a, 16'h838b, 16'h7b6a, 16'h20e3, 16'h62a9, 16'h62ea, 16'h39c8, 16'h31a7, 16'h524a, 16'hb513, 16'hc594, 16'hc554, 16'hb512, 16'hacd1, 16'hacb1, 16'ha490, 16'h9c4f, 16'h93ee, 16'h7b2b, 16'h8bcd, 16'h836c, 16'h7b2b, 16'h6aa9, 16'h6268, 16'h5227, 16'h526, 16'h5227, 16'h73a, 16'h5227, 16'h527, 16'h49e6, 16'h5a68, 16'h4184, 16'h3964, 16'h3185, 16'h841, 16'h840, 16'h20e2, 16'h3984, 16'h49e5, 16'h5a46, 16'h49c5, 16'h49c5, 16'h49e6, 16'h6289, 16'h6289, 16'h5227, 16'h41c5, 16'h4a6, 16'h4184, 16'h3984, 16'h3984, 16'h3963, 16'h3122, 16'h3143, 16'h3143, 16'h18c2, 16'h840, 16'h840, 16'h861, 16'h1061, 16'h1081, 16'h1081, 16'h18c2, 16'h20e2, 16'h18a1, 16'h18c2, 16'h212, 16'h212, 16'h20e2, 16'h20e2, 16'h20e3, 16'h20e2, 16'h18c2, 16'h18a2, 16'h18c2, 16'h20c3, 16'h7b2c, 16'hde16, 16'hde36, 16'hde36, 16'hde16, 16'hde16, 16'hde16, 16'hd616, 16'hd616, 16'hd616, 16'hd5f6, 16'hd5f6, 16'hd5f5, 16'hd5d5, 16'hd5d5, 16'hd5d5, 16'hd5d5, 16'hd5d5, 16'hd5b5, 16'hcdb5, 16'hcdb5, 16'hcdb5, 16'hcdb4, 16'hcdb4, 16'hcd94, 16'hcd94, 16'hcd94, 16'hc594, 16'hc594, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc553, 16'hc553, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd32, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd33, 16'ha450, 16'h3165, 16'h20e3, 16'h20e2, 16'h20c2, 16'h18c2, 16'h1061, 16'h020, 16'h020, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h7bab, 16'h83cc, 16'h8bec, 16'h8cd, 16'h8c2d, 16'h942d, 16'h944e, 16'h944f, 16'h9c6f, 16'h9c6f, 16'h9c6f, 16'h9c8f, 16'h9c8f, 16'h9c8f, 16'h9c8f, 16'h9c8f, 16'h9c6e, 16'h734a, 16'h18c2, 16'h860, 16'h860, 16'h1081, 16'h4a7, 16'h3164, 16'h1081, 16'h1081, 16'h18a1, 16'h10a1, 16'h10c1, 16'h1081, 16'h1081, 16'h881, 16'h1082, 16'h293, 16'h5226, 16'h5a68, 16'h62a9, 16'h732a, 16'h7329, 16'h20e3, 16'h6289, 16'h5aaa, 16'h31c8, 16'h31a8, 16'h62ab, 16'hbd53, 16'hc574, 16'hc553, 16'hb512, 16'hacd1, 16'hacb0, 16'ha490, 16'h9c6f, 16'h94e, 16'h7b2b, 16'h8bad, 16'h836c, 16'h7ba, 16'h6aa9, 16'h6268, 16'h5a68, 16'h5227, 16'h5227, 16'h73a, 16'h5227, 16'h527, 16'h526, 16'h5a68, 16'h4184, 16'h3984, 16'h39a5, 16'h861, 16'h020, 16'h18c2, 16'h293, 16'h3143, 16'h3963, 16'h3964, 16'h41a5, 16'h5a27, 16'h6ac9, 16'h6289, 16'h5227, 16'h41c5, 16'h4a6, 16'h41a4, 16'h3984, 16'h3983, 16'h3963, 16'h3143, 16'h3143, 16'h3963, 16'h20c2, 16'h820, 16'h020, 16'h020, 16'h020, 16'h820, 16'h820, 16'h820, 16'h18a2, 16'h18a1, 16'h1040, 16'h1081, 16'h18c2, 16'h18c2, 16'h18c2, 16'h18a2, 16'h1062, 16'h840, 16'h840, 16'h840, 16'h1061, 16'h73b, 16'hde36, 16'hde37, 16'hde36, 16'hde36, 16'hde36, 16'hde16, 16'hde16, 16'hd616, 16'hd616, 16'hd616, 16'hd5f6, 16'hd5f6, 16'hd5f5, 16'hd5d5, 16'hd5d5, 16'hd5d5, 16'hd5b5, 16'hd5b5, 16'hd5b5, 16'hcdb5, 16'hcdb5, 16'hcdb5, 16'hcdb4, 16'hcd94, 16'hcd94, 16'hcd94, 16'hc594, 16'hc594, 16'hc574, 16'hc574, 16'hc574, 16'hc573, 16'hc574, 16'hc553, 16'hc553, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd32, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd33, 16'h9c4f, 16'h3165, 16'h20e3, 16'h20e2, 16'h18e2, 16'h18c2, 16'h1061, 16'h020, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h83ec, 16'h8cd, 16'h8cd, 16'h942d, 16'h944e, 16'h946f, 16'h9c6f, 16'h9c8f, 16'h9c8f, 16'h9c8f, 16'h9c8f, 16'ha4af, 16'h9caf, 16'h9caf, 16'h9c8f, 16'h9c8f, 16'h9c8f, 16'h7b8b, 16'h3985, 16'h213, 16'h18c2, 16'h18a2, 16'h4a27, 16'h41e6, 16'h1081, 16'h1081, 16'h1060, 16'h861, 16'h861, 16'h861, 16'h861, 16'h861, 16'h1061, 16'h1081, 16'h1881, 16'h18a2, 16'h18c2, 16'h2123, 16'h3163, 16'h18a2, 16'h62a9, 16'h5a8a, 16'h31c8, 16'h31a8, 16'h6aec, 16'hc554, 16'hc574, 16'hc573, 16'hb532, 16'hacd1, 16'hacb1, 16'ha490, 16'h9c6f, 16'h94e, 16'h73b, 16'h8bcd, 16'h836c, 16'h7bb, 16'h6aca, 16'h6288, 16'h5a48, 16'h527, 16'h5228, 16'h73b, 16'h5227, 16'h527, 16'h49e6, 16'h5a68, 16'h3964, 16'h3964, 16'h41c6, 16'h861, 16'h820, 16'h2923, 16'h41a4, 16'h41a4, 16'h49c5, 16'h49c5, 16'h51e6, 16'h5a48, 16'h6ac9, 16'h62a9, 16'h5227, 16'h41c6, 16'h4a6, 16'h41a4, 16'h3984, 16'h3983, 16'h3963, 16'h3964, 16'h3963, 16'h3963, 16'h20c2, 16'h820, 16'h820, 16'h020, 16'h020, 16'h840, 16'h840, 16'h1060, 16'h1081, 16'h18a1, 16'h1081, 16'h840, 16'h841, 16'h1061, 16'h1081, 16'h1082, 16'h861, 16'h840, 16'h040, 16'h840, 16'h1061, 16'h73c, 16'hde36, 16'hde37, 16'hde36, 16'hde36, 16'hde36, 16'hde16, 16'hde16, 16'hd616, 16'hde16, 16'hd616, 16'hd5f6, 16'hd5f6, 16'hd5f5, 16'hd5f5, 16'hd5d5, 16'hd5d5, 16'hd5d5, 16'hd5d5, 16'hd5d5, 16'hcdb5, 16'hcdb5, 16'hcdb5, 16'hcdb5, 16'hcd94, 16'hcd94, 16'hcd94, 16'hc594, 16'hc594, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc553, 16'hc553, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd33, 16'hbd13, 16'h9cf, 16'h3145, 16'h20e2, 16'h20e2, 16'h20e2, 16'h18c2, 16'h1061, 16'h020, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h8cd, 16'h942e, 16'h944e, 16'h9c6e, 16'h9c8f, 16'h9c8f, 16'ha4b0, 16'ha4b0, 16'ha4b0, 16'ha4b0, 16'ha4b0, 16'ha4b0, 16'ha4b0, 16'ha4af, 16'ha4af, 16'h9c8f, 16'h9c8f, 16'h9c8f, 16'h942e, 16'h8bed, 16'h7b8c, 16'h732b, 16'h6ae9, 16'h4a27, 16'h1081, 16'h1061, 16'h1080, 16'h880, 16'h860, 16'h860, 16'h860, 16'h860, 16'h860, 16'h860, 16'h860, 16'h840, 16'h861, 16'h861, 16'h10a1, 16'h18c2, 16'h6289, 16'h528a, 16'h39c8, 16'h3188, 16'h732d, 16'hc574, 16'hc574, 16'hc573, 16'hbd32, 16'hb4f1, 16'hacb1, 16'ha4b0, 16'ha470, 16'h94e, 16'h73b, 16'h8bcd, 16'h838c, 16'h7b2b, 16'h6aa9, 16'h6268, 16'h5a48, 16'h5227, 16'h5227, 16'h73b, 16'h5227, 16'h527, 16'h527, 16'h6268, 16'h41a4, 16'h41a5, 16'h49e7, 16'h861, 16'h840, 16'h2923, 16'h49c4, 16'h41a4, 16'h4184, 16'h4184, 16'h49e5, 16'h5a47, 16'h6aca, 16'h62a9, 16'h5227, 16'h41c6, 16'h4a6, 16'h41a4, 16'h39a4, 16'h3983, 16'h3963, 16'h3963, 16'h3963, 16'h3963, 16'h20c2, 16'h820, 16'h020, 16'h020, 16'h840, 16'h1081, 16'h1061, 16'h1081, 16'h1061, 16'h1061, 16'h18a1, 16'h861, 16'h020, 16'h020, 16'h040, 16'h841, 16'h840, 16'h040, 16'h040, 16'h840, 16'h1061, 16'h73b, 16'hde37, 16'hde37, 16'hde37, 16'hde36, 16'hde36, 16'hde36, 16'hde16, 16'hde16, 16'hde16, 16'hd616, 16'hd616, 16'hd5f6, 16'hd5f6, 16'hd5f6, 16'hd5f5, 16'hd5d5, 16'hd5d5, 16'hd5d5, 16'hd5d5, 16'hcdd5, 16'hcdb5, 16'hcdb5, 16'hcdb5, 16'hcdb5, 16'hcd94, 16'hcd94, 16'hcd94, 16'hc594, 16'hc594, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc573, 16'hc553, 16'hc553, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hbd12, 16'hbd12, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd13, 16'hbd13, 16'h94f, 16'h3144, 16'h20e2, 16'h20c2, 16'h20e2, 16'h20c2, 16'h1061, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h944e, 16'h9c6f, 16'h9c8f, 16'h9c8f, 16'ha4b0, 16'ha4b0, 16'ha4d0, 16'ha4d0, 16'ha4d0, 16'ha4d0, 16'ha4d0, 16'ha4d0, 16'ha4d0, 16'ha4b0, 16'ha4b0, 16'ha4af, 16'h9caf, 16'h9c90, 16'h9c6f, 16'h9c6f, 16'h946f, 16'h942e, 16'h732a, 16'h4a26, 16'h10a1, 16'h1061, 16'h1060, 16'h1061, 16'h1061, 16'h1060, 16'h860, 16'h860, 16'h861, 16'h860, 16'h840, 16'h020, 16'h020, 16'h820, 16'h840, 16'h10a1, 16'h5a88, 16'h526a, 16'h39c8, 16'h31a8, 16'h734d, 16'hbd53, 16'hc574, 16'hc574, 16'hb512, 16'hb4d2, 16'hacb1, 16'ha4b0, 16'ha470, 16'h94e, 16'h7b2b, 16'h93ce, 16'h8b8d, 16'h7b4c, 16'h6aa9, 16'h5a48, 16'h5a28, 16'h5227, 16'h5248, 16'h732b, 16'h5227, 16'h527, 16'h49e6, 16'h6288, 16'h41a4, 16'h4184, 16'h4a7, 16'h861, 16'h840, 16'h293, 16'h4184, 16'h3123, 16'h3964, 16'h41a4, 16'h49c5, 16'h6268, 16'h72ca, 16'h6aa9, 16'h5227, 16'h41c5, 16'h4a6, 16'h41a4, 16'h3984, 16'h3984, 16'h3963, 16'h3963, 16'h3963, 16'h3964, 16'h20e2, 16'h840, 16'h020, 16'h020, 16'h1081, 16'h10a1, 16'h1060, 16'h1080, 16'h1060, 16'h1061, 16'h1081, 16'h10a1, 16'h020, 16'h020, 16'h020, 16'h040, 16'h040, 16'h040, 16'h040, 16'h840, 16'h1062, 16'h73b, 16'hde37, 16'hde37, 16'hde37, 16'hde37, 16'hde36, 16'hde36, 16'hde36, 16'hde16, 16'hde16, 16'hd616, 16'hd616, 16'hd5f6, 16'hd5f6, 16'hd5f6, 16'hd5f5, 16'hd5d5, 16'hd5d5, 16'hd5d5, 16'hd5d5, 16'hcdd5, 16'hcdd5, 16'hcdb5, 16'hcdb5, 16'hcdb5, 16'hcdb4, 16'hcd94, 16'hcd94, 16'hc594, 16'hc594, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc553, 16'hc553, 16'hc553, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hbd32, 16'hbd12, 16'hbd12, 16'hbd12, 16'hb512, 16'hbd12, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd32, 16'hbd12, 16'hbd33, 16'hbd12, 16'h93ee, 16'h3145, 16'h20e3, 16'h20c2, 16'h20c2, 16'h20c2, 16'h1061, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h9c8f, 16'h9cb0, 16'ha4b0, 16'ha4d0, 16'ha4d0, 16'ha4d0, 16'hacd0, 16'hacf0, 16'ha4f0, 16'ha4d0, 16'ha4d0, 16'ha4d0, 16'ha4d0, 16'ha4b0, 16'ha4b0, 16'ha4af, 16'h9caf, 16'h9c8f, 16'h9c6f, 16'h946f, 16'h944e, 16'h942d, 16'h6ba, 16'h49e6, 16'h10a1, 16'h1061, 16'h1061, 16'h1081, 16'h1061, 16'h1060, 16'h860, 16'h860, 16'h860, 16'h860, 16'h860, 16'h040, 16'h840, 16'h860, 16'h841, 16'h1061, 16'h5268, 16'h526a, 16'h39c8, 16'h31a8, 16'h734d, 16'hbd53, 16'hc574, 16'hc574, 16'hbd32, 16'hb4f2, 16'hacd1, 16'hacb0, 16'ha470, 16'h94e, 16'h7b2b, 16'h93ee, 16'h8bad, 16'h7b4b, 16'h6aa9, 16'h5a48, 16'h5228, 16'h5a28, 16'h5a48, 16'h732a, 16'h5247, 16'h49e6, 16'h41a5, 16'h5a68, 16'h41a4, 16'h4185, 16'h5248, 16'h1081, 16'h840, 16'h2923, 16'h49e5, 16'h49a5, 16'h49a5, 16'h49c5, 16'h49c5, 16'h5a68, 16'h72ea, 16'h6aa9, 16'h5227, 16'h49e6, 16'h4a6, 16'h39a4, 16'h3984, 16'h3984, 16'h3983, 16'h3963, 16'h3164, 16'h3964, 16'h20e2, 16'h840, 16'h040, 16'h1081, 16'h18a2, 16'h860, 16'h860, 16'h1081, 16'h1061, 16'h860, 16'h860, 16'h18c2, 16'h841, 16'h020, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h841, 16'h1062, 16'h73c, 16'hde37, 16'hde37, 16'hde37, 16'hde37, 16'hde37, 16'hde36, 16'hde36, 16'hde16, 16'hde16, 16'hd616, 16'hd5f6, 16'hd5f6, 16'hd5f6, 16'hd5f6, 16'hd5f5, 16'hd5d5, 16'hd5d5, 16'hd5d5, 16'hd5d5, 16'hcdd5, 16'hcdd5, 16'hcdb5, 16'hcdb5, 16'hcdb5, 16'hcdb4, 16'hcd94, 16'hcd94, 16'hc594, 16'hc594, 16'hc594, 16'hc574, 16'hc574, 16'hc574, 16'hc573, 16'hc553, 16'hc553, 16'hc553, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hbd32, 16'hbd12, 16'hbd12, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hb512, 16'h8bce, 16'h3144, 16'h20e2, 16'h20e2, 16'h20c2, 16'h20c2, 16'h1061, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'ha4af, 16'h9c8f, 16'ha4b0, 16'ha4b0, 16'ha4b0, 16'h9c6f, 16'hacf1, 16'ha4d1, 16'ha4d0, 16'hacf1, 16'hacf0, 16'ha4d0, 16'ha4d0, 16'ha4d0, 16'ha4b0, 16'ha4af, 16'h9c8f, 16'h9c6f, 16'h9c6f, 16'h944f, 16'h944e, 16'h942d, 16'h6ba, 16'h49e6, 16'h10a1, 16'h1081, 16'h1081, 16'h1081, 16'h1081, 16'h1060, 16'h860, 16'h860, 16'h860, 16'h860, 16'h860, 16'h840, 16'h861, 16'h1081, 16'h1081, 16'h1062, 16'h5a68, 16'h5a8a, 16'h39c9, 16'h39a8, 16'h73c, 16'hb533, 16'hc574, 16'hc574, 16'hbd33, 16'hb4f2, 16'hacd1, 16'hacb1, 16'ha470, 16'h94e, 16'h7b2b, 16'h93ee, 16'h8bad, 16'h836c, 16'h6aa9, 16'h5a27, 16'h5228, 16'h5a48, 16'h5247, 16'h732b, 16'h5227, 16'h4a7, 16'h49e7, 16'h5a89, 16'h41a5, 16'h49a5, 16'h5a88, 16'h18a2, 16'h840, 16'h3143, 16'h5a46, 16'h5a25, 16'h5a5, 16'h51e4, 16'h5a25, 16'h5a67, 16'h73a, 16'h6aea, 16'h5247, 16'h41a5, 16'h4a6, 16'h41a4, 16'h3984, 16'h3984, 16'h3983, 16'h3964, 16'h3964, 16'h3983, 16'h20e2, 16'h840, 16'h840, 16'h861, 16'h840, 16'h840, 16'h840, 16'h1081, 16'h1081, 16'h860, 16'h860, 16'h10a1, 16'h1081, 16'h020, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h841, 16'h1062, 16'h73c, 16'hde37, 16'hde37, 16'hde37, 16'hde37, 16'hde37, 16'hde36, 16'hde16, 16'hde16, 16'hde16, 16'hd616, 16'hd5f6, 16'hd5f6, 16'hd5f6, 16'hd5f6, 16'hd5f5, 16'hd5d5, 16'hd5d5, 16'hd5d5, 16'hd5d5, 16'hd5d5, 16'hcdd5, 16'hcdb5, 16'hcdb5, 16'hcdb5, 16'hcdb4, 16'hcd94, 16'hcd94, 16'hcd94, 16'hc594, 16'hc594, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc573, 16'hc553, 16'hc553, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hbd12, 16'hbd12, 16'hb512, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb512, 16'hb512, 16'hb4f2, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hbd12, 16'hbd12, 16'hb512, 16'hb512, 16'hb4f2, 16'h8bad, 16'h3144, 16'h20e2, 16'h20e2, 16'h20e2, 16'h20c2, 16'h1061, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'ha4d0, 16'h9c8f, 16'ha4b0, 16'ha4b0, 16'ha4d1, 16'ha4b0, 16'hacf1, 16'hacf1, 16'ha4d0, 16'ha4b0, 16'hacf1, 16'ha4d1, 16'ha4d0, 16'ha4d0, 16'ha4b0, 16'h9caf, 16'h9c8f, 16'h9c6f, 16'h9c6f, 16'h944f, 16'h944e, 16'h942d, 16'h6ba, 16'h41e6, 16'h10a1, 16'h1081, 16'h861, 16'h1061, 16'h1081, 16'h1080, 16'h860, 16'h860, 16'h860, 16'h860, 16'h840, 16'h840, 16'h840, 16'h18c2, 16'h2924, 16'h1082, 16'h5a68, 16'h62cb, 16'h39e9, 16'h31c8, 16'h62cb, 16'hacd2, 16'hbd53, 16'hc574, 16'hbd53, 16'hacf2, 16'hacb1, 16'ha490, 16'ha470, 16'h94e, 16'h7b4b, 16'h93ee, 16'h8bad, 16'h836c, 16'h6289, 16'h5227, 16'h527, 16'h5248, 16'h4a7, 16'h732b, 16'h5227, 16'h4a7, 16'h4a7, 16'h62a9, 16'h41a5, 16'h4184, 16'h62a9, 16'h20c3, 16'h840, 16'h41a5, 16'h5a67, 16'h51e5, 16'h5a26, 16'h526, 16'h526, 16'h527, 16'h6ae9, 16'h6aea, 16'h5247, 16'h41a5, 16'h5226, 16'h41a4, 16'h3984, 16'h3984, 16'h3983, 16'h3984, 16'h3983, 16'h3983, 16'h212, 16'h840, 16'h840, 16'h020, 16'h020, 16'h020, 16'h840, 16'h1081, 16'h1081, 16'h860, 16'h860, 16'h861, 16'h1081, 16'h020, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h841, 16'h1062, 16'h732b, 16'hde37, 16'hde37, 16'hde37, 16'hde37, 16'hde37, 16'hde36, 16'hde16, 16'hde16, 16'hde16, 16'hd616, 16'hd616, 16'hd5f6, 16'hd5f6, 16'hd5f5, 16'hd5f5, 16'hd5d5, 16'hd5d5, 16'hd5d5, 16'hd5d5, 16'hd5d5, 16'hcdd5, 16'hcdb5, 16'hcdb5, 16'hcdb5, 16'hcdb4, 16'hcd94, 16'hcd94, 16'hcd94, 16'hc594, 16'hc594, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc573, 16'hc553, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hbd12, 16'hb512, 16'hbd12, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb512, 16'hb512, 16'hb4f2, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'h83ad, 16'h3144, 16'h20e2, 16'h20c2, 16'h20c2, 16'h20c2, 16'h1061, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'had11, 16'hacf1, 16'had12, 16'had11, 16'had11, 16'had11, 16'had11, 16'hacf1, 16'ha4d0, 16'ha490, 16'ha4f1, 16'ha4d1, 16'ha4d0, 16'ha4d0, 16'h9cb0, 16'h9c8f, 16'h9c8f, 16'h9c6f, 16'h9c6f, 16'h944f, 16'h944e, 16'h942e, 16'h6ba, 16'h41e6, 16'h10a1, 16'h861, 16'h860, 16'h860, 16'h1080, 16'h1061, 16'h1061, 16'h861, 16'h860, 16'h860, 16'h860, 16'h18c2, 16'h10a2, 16'h18e2, 16'h2943, 16'h1082, 16'h5a68, 16'h734c, 16'h3a9, 16'h31c8, 16'h526a, 16'ha471, 16'hb512, 16'hc574, 16'hbd33, 16'hb4f2, 16'hacb1, 16'ha490, 16'h9c70, 16'h94e, 16'h7b4c, 16'h93ee, 16'h8bcd, 16'h836c, 16'h6268, 16'h5227, 16'h527, 16'h5248, 16'h49e6, 16'h732b, 16'h5228, 16'h527, 16'h527, 16'h62a9, 16'h49c5, 16'h41a5, 16'h6bb, 16'h3985, 16'h840, 16'h2923, 16'h49c5, 16'h49a4, 16'h49a4, 16'h49a4, 16'h49a4, 16'h49c5, 16'h527, 16'h5228, 16'h5a28, 16'h5227, 16'h5227, 16'h4184, 16'h3984, 16'h3984, 16'h3984, 16'h3984, 16'h3984, 16'h3984, 16'h212, 16'h840, 16'h840, 16'h020, 16'h020, 16'h020, 16'h840, 16'h1081, 16'h1081, 16'h1060, 16'h1061, 16'h10a1, 16'h861, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h041, 16'h841, 16'h862, 16'h73c, 16'hde37, 16'hde37, 16'hde37, 16'hde37, 16'hde37, 16'hde36, 16'hde16, 16'hde16, 16'hde16, 16'hd616, 16'hd5f6, 16'hd5f6, 16'hd5f6, 16'hd5f5, 16'hd5f5, 16'hd5d5, 16'hd5d5, 16'hd5d5, 16'hd5d5, 16'hd5d5, 16'hd5d5, 16'hcdb5, 16'hcdb5, 16'hcdb5, 16'hcdb4, 16'hcd94, 16'hcd94, 16'hc594, 16'hc594, 16'hc574, 16'hc574, 16'hc574, 16'hc573, 16'hc573, 16'hc573, 16'hc553, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'h83ac, 16'h3144, 16'h20e2, 16'h20c2, 16'h20c2, 16'h18c2, 16'h1061, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'had11, 16'hacd1, 16'had12, 16'had11, 16'had11, 16'had11, 16'hacf1, 16'hacf1, 16'ha4d0, 16'ha4b0, 16'ha4d1, 16'ha4d1, 16'ha4d0, 16'ha4d0, 16'ha4b0, 16'h9cb0, 16'h9c90, 16'h9c8f, 16'h9c6f, 16'h946f, 16'h944f, 16'h942e, 16'h6ba, 16'h39c5, 16'h10a1, 16'h861, 16'h860, 16'h1061, 16'h1061, 16'h1060, 16'h860, 16'h861, 16'h860, 16'h860, 16'h1081, 16'h39a5, 16'h2964, 16'h1061, 16'h1081, 16'h1061, 16'h5a68, 16'h83ad, 16'h4229, 16'h31a8, 16'h39c8, 16'h838d, 16'h9c50, 16'hbd33, 16'hbd33, 16'hb512, 16'hacd1, 16'ha490, 16'h9c4f, 16'h93ee, 16'h834c, 16'h94e, 16'h8bcd, 16'h7b4b, 16'h5a68, 16'h527, 16'h4a7, 16'h5227, 16'h41c6, 16'h7b2b, 16'h5248, 16'h5227, 16'h4a7, 16'h6289, 16'h49e6, 16'h3164, 16'h3984, 16'h18a2, 16'h840, 16'h18c2, 16'h41c6, 16'h5227, 16'h5227, 16'h527, 16'h49e6, 16'h49e6, 16'h5248, 16'h6aaa, 16'h5a28, 16'h49c6, 16'h41c6, 16'h3984, 16'h3984, 16'h3984, 16'h3984, 16'h3984, 16'h3984, 16'h39a4, 16'h212, 16'h840, 16'h840, 16'h840, 16'h020, 16'h020, 16'h840, 16'h1081, 16'h1081, 16'h1081, 16'h10a1, 16'h1081, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h041, 16'h041, 16'h841, 16'h1062, 16'h73c, 16'hde37, 16'hde57, 16'hde37, 16'hde37, 16'hde37, 16'hde16, 16'hde16, 16'hde16, 16'hde16, 16'hd616, 16'hd5f6, 16'hd5f6, 16'hd5f6, 16'hd5f6, 16'hd5f5, 16'hd5d5, 16'hd5d5, 16'hd5d5, 16'hd5d5, 16'hd5d5, 16'hcdb5, 16'hcdb5, 16'hcdb5, 16'hcdb4, 16'hcdb4, 16'hcdb4, 16'hcd94, 16'hc594, 16'hc594, 16'hc574, 16'hc574, 16'hc573, 16'hc573, 16'hc573, 16'hc553, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'h838c, 16'h2944, 16'h20e2, 16'h20e2, 16'h20c2, 16'h18c2, 16'h1061, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'hb531, 16'hacf1, 16'hb532, 16'hb532, 16'had12, 16'had11, 16'hacf1, 16'hacf1, 16'ha4d0, 16'ha4b0, 16'ha4f0, 16'ha4d0, 16'ha4d0, 16'ha4d0, 16'ha4b0, 16'h9cb0, 16'h9c90, 16'h9c90, 16'h9c6f, 16'h9c6f, 16'h944f, 16'h944e, 16'h6ba, 16'h39a5, 16'h10a1, 16'h861, 16'h860, 16'h861, 16'h881, 16'h1061, 16'h861, 16'h861, 16'h860, 16'h860, 16'h860, 16'h10a2, 16'h10a1, 16'h840, 16'h840, 16'h841, 16'h5247, 16'h94d, 16'h62cb, 16'h3188, 16'h3187, 16'h6aeb, 16'h8b8d, 16'hacb1, 16'hb533, 16'hb533, 16'hb4f2, 16'ha4b1, 16'h9c4f, 16'h8bcd, 16'h836c, 16'h94e, 16'h93cd, 16'h7b2b, 16'h5a48, 16'h4a7, 16'h49e7, 16'h49e7, 16'h3985, 16'h7b4b, 16'h5a68, 16'h4a6, 16'h49e6, 16'h5a68, 16'h49e5, 16'h3163, 16'h20e2, 16'h861, 16'h820, 16'h10a2, 16'h49e6, 16'h5a68, 16'h5227, 16'h5a48, 16'h6288, 16'h6ac9, 16'h7b2b, 16'h73a, 16'h5227, 16'h49e6, 16'h4a6, 16'h3984, 16'h3984, 16'h3984, 16'h3984, 16'h41a4, 16'h41a4, 16'h41a4, 16'h2923, 16'h1081, 16'h881, 16'h861, 16'h820, 16'h020, 16'h840, 16'h1061, 16'h1081, 16'h1081, 16'h1081, 16'h860, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h041, 16'h041, 16'h861, 16'h1062, 16'h73c, 16'hde37, 16'hde57, 16'hde37, 16'hde36, 16'hde36, 16'hde16, 16'hde16, 16'hde16, 16'hd616, 16'hd616, 16'hd5f6, 16'hd5f6, 16'hd5f6, 16'hd5f5, 16'hd5d5, 16'hd5d5, 16'hd5d5, 16'hd5d5, 16'hd5d5, 16'hd5d5, 16'hcdb5, 16'hcdb5, 16'hcdb4, 16'hcdb4, 16'hcdb4, 16'hcd94, 16'hc594, 16'hc594, 16'hc594, 16'hc574, 16'hc574, 16'hc574, 16'hc573, 16'hc553, 16'hc553, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hb512, 16'hbd12, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4d1, 16'h7b6c, 16'h2924, 16'h20e2, 16'h20e2, 16'h20c2, 16'h18c2, 16'h1061, 16'h020, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'hb552, 16'hb532, 16'hb552, 16'hb552, 16'hb552, 16'hb532, 16'hb532, 16'had11, 16'hacf1, 16'ha4f1, 16'hacf1, 16'ha4d1, 16'ha4d0, 16'ha4d0, 16'ha4b0, 16'ha4b0, 16'h9cb0, 16'h9c90, 16'h9c8f, 16'h9c6f, 16'h946f, 16'h944e, 16'h6ba, 16'h39a5, 16'h10a1, 16'h861, 16'h860, 16'h1061, 16'h1081, 16'h1061, 16'h1061, 16'h861, 16'h860, 16'h860, 16'h860, 16'h040, 16'h840, 16'h861, 16'h10a2, 16'h1082, 16'h5248, 16'h942d, 16'h8bed, 16'h62aa, 16'h39c7, 16'h5a49, 16'h836d, 16'h942f, 16'hb4f2, 16'hb512, 16'hb512, 16'hacb1, 16'ha470, 16'h8bad, 16'h834c, 16'h93ed, 16'h8bcd, 16'h7b2b, 16'h5a48, 16'h49e7, 16'h49e6, 16'h3985, 16'h3965, 16'h7b4b, 16'h6288, 16'h3985, 16'h3985, 16'h4a7, 16'h49e5, 16'h3123, 16'h20e2, 16'h18a2, 16'h1061, 16'h861, 16'h49e6, 16'h6aa9, 16'h5a47, 16'h5a68, 16'h6ac9, 16'h72ea, 16'h836c, 16'h73a, 16'h5227, 16'h41a5, 16'h49e6, 16'h3984, 16'h41a4, 16'h41a4, 16'h41a4, 16'h41a4, 16'h41a4, 16'h41a4, 16'h292, 16'h860, 16'h840, 16'h840, 16'h00, 16'h00, 16'h820, 16'h1061, 16'h18a1, 16'h1081, 16'h1081, 16'h860, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h841, 16'h841, 16'h1062, 16'h73c, 16'hde37, 16'hde37, 16'hde36, 16'hde36, 16'hde16, 16'hde16, 16'hde16, 16'hd616, 16'hd616, 16'hd5f6, 16'hd5f6, 16'hd5f6, 16'hd5f6, 16'hd5d5, 16'hd5d5, 16'hd5d5, 16'hd5d5, 16'hd5d5, 16'hd5d5, 16'hd5b5, 16'hcdb5, 16'hcdb5, 16'hcdb4, 16'hcdb4, 16'hcd94, 16'hcd94, 16'hc594, 16'hc594, 16'hc574, 16'hc574, 16'hc574, 16'hc573, 16'hc573, 16'hc573, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd32, 16'hbd12, 16'hbd12, 16'hbd32, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hacd1, 16'h7b4c, 16'h2924, 16'h20e2, 16'h20e2, 16'h20c2, 16'h20c2, 16'h1061, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'hb552, 16'hb552, 16'hb552, 16'hb532, 16'hb532, 16'hb532, 16'had32, 16'had12, 16'had11, 16'hacf1, 16'hacf1, 16'ha4f1, 16'ha4d0, 16'ha4d0, 16'ha4d0, 16'ha4b0, 16'ha4b0, 16'h9c90, 16'h9c8f, 16'h9c6f, 16'h946f, 16'h944e, 16'h6b2a, 16'h31a4, 16'h10a1, 16'h861, 16'h860, 16'h1060, 16'h1061, 16'h1061, 16'h1061, 16'h860, 16'h860, 16'h860, 16'h840, 16'h040, 16'h840, 16'h861, 16'h18e3, 16'h18c3, 16'h5247, 16'h942d, 16'h942e, 16'h942e, 16'h8bcd, 16'h838c, 16'h8bcd, 16'h8bad, 16'ha4b0, 16'hacd1, 16'hb512, 16'hacd2, 16'ha470, 16'h838c, 16'h836c, 16'h93ee, 16'h8b8d, 16'h72ea, 16'h5a48, 16'h49e6, 16'h41a5, 16'h2923, 16'h3165, 16'h7b4b, 16'h62a9, 16'h3164, 16'h3985, 16'h3984, 16'h3164, 16'h3123, 16'h293, 16'h213, 16'h18a2, 16'h020, 16'h293, 16'h6288, 16'h5a68, 16'h6ac9, 16'h6ac9, 16'h49c6, 16'h5a47, 16'h5a48, 16'h5247, 16'h3985, 16'h41c6, 16'h41a4, 16'h41a4, 16'h41a4, 16'h41a4, 16'h3984, 16'h41a4, 16'h41a4, 16'h212, 16'h840, 16'h840, 16'h820, 16'h00, 16'h00, 16'h020, 16'h1061, 16'h18a1, 16'h1081, 16'h1081, 16'h860, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h840, 16'h841, 16'h1062, 16'h73c, 16'hde37, 16'hde37, 16'hde36, 16'hde36, 16'hde16, 16'hde16, 16'hd616, 16'hd616, 16'hd5f6, 16'hd5f6, 16'hd5f6, 16'hd5f5, 16'hd5f5, 16'hd5f5, 16'hd5d5, 16'hd5d5, 16'hcdd5, 16'hcdb5, 16'hcdb5, 16'hcdb5, 16'hcdb5, 16'hcdb5, 16'hcdb4, 16'hcd94, 16'hcd94, 16'hcd94, 16'hc594, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc573, 16'hc553, 16'hc553, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4d2, 16'hb4f2, 16'hb4f1, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hacd1, 16'h7b4c, 16'h2924, 16'h20e2, 16'h20e2, 16'h20c2, 16'h18c2, 16'h1061, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'hb552, 16'hb552, 16'hb552, 16'hb552, 16'hb532, 16'hb532, 16'had32, 16'had12, 16'had11, 16'had11, 16'hacf1, 16'ha4f1, 16'ha4f1, 16'ha4d0, 16'ha4d0, 16'ha4d0, 16'ha4b0, 16'h9cb0, 16'h9c90, 16'h942e, 16'h83ac, 16'h83ac, 16'h6b9, 16'h3164, 16'h1081, 16'h861, 16'h861, 16'h861, 16'h1061, 16'h1061, 16'h1060, 16'h860, 16'h861, 16'h860, 16'h860, 16'h040, 16'h040, 16'h881, 16'h1081, 16'h861, 16'h5227, 16'h942d, 16'h942e, 16'h942d, 16'h942e, 16'h9c6f, 16'h94e, 16'h838c, 16'h942f, 16'ha490, 16'hacd1, 16'hb4f2, 16'ha490, 16'h7b4b, 16'h7b4b, 16'h8bad, 16'h7b4c, 16'h73a, 16'h6288, 16'h49e6, 16'h3985, 16'h20c2, 16'h3165, 16'h7b4b, 16'h62a9, 16'h3964, 16'h3985, 16'h293, 16'h293, 16'h3144, 16'h293, 16'h2924, 16'h20c3, 16'h820, 16'h820, 16'h3164, 16'h5247, 16'h5a88, 16'h49e6, 16'h3144, 16'h41a5, 16'h5227, 16'h5a68, 16'h3124, 16'h41a5, 16'h41a5, 16'h41c5, 16'h41c5, 16'h41a4, 16'h3984, 16'h4184, 16'h41a4, 16'h212, 16'h840, 16'h840, 16'h820, 16'h00, 16'h00, 16'h020, 16'h1061, 16'h18a1, 16'h1081, 16'h1081, 16'h1061, 16'h840, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h041, 16'h841, 16'h1062, 16'h73b, 16'hde36, 16'hde36, 16'hde16, 16'hde16, 16'hde16, 16'hd616, 16'hd616, 16'hd5f6, 16'hd5f6, 16'hd5f6, 16'hd5f5, 16'hd5f5, 16'hd5d5, 16'hd5d5, 16'hd5d5, 16'hcdd5, 16'hcdb5, 16'hcdb5, 16'hcdb5, 16'hcdb5, 16'hcdb5, 16'hcdb4, 16'hcd94, 16'hcd94, 16'hcd94, 16'hc594, 16'hc574, 16'hc574, 16'hc574, 16'hc573, 16'hc573, 16'hc573, 16'hc553, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4f1, 16'hb4f1, 16'hb4f2, 16'hb4d1, 16'hb4d1, 16'hb4f1, 16'hb4d1, 16'hb4d2, 16'hb4d2, 16'hb4d1, 16'hacb1, 16'h7b4b, 16'h2924, 16'h20e2, 16'h20c2, 16'h18c2, 16'h18c2, 16'h1061, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'hb552, 16'hb552, 16'hb552, 16'hb552, 16'hb552, 16'hb532, 16'hb532, 16'had32, 16'had11, 16'had11, 16'hacf1, 16'hacf1, 16'ha4f1, 16'ha4d1, 16'ha4d0, 16'ha4d0, 16'ha4b0, 16'h9cb0, 16'h9c90, 16'h734b, 16'h2923, 16'h2923, 16'h39c5, 16'h2923, 16'h1081, 16'h861, 16'h861, 16'h861, 16'h861, 16'h1061, 16'h861, 16'h861, 16'h861, 16'h860, 16'h860, 16'h840, 16'h840, 16'h860, 16'h840, 16'h841, 16'h4a27, 16'h94e, 16'h942e, 16'h942e, 16'h942e, 16'h9c6f, 16'h9c2d, 16'h8bac, 16'h93ee, 16'h9c4f, 16'ha470, 16'hacb1, 16'ha4b0, 16'h73a, 16'h49c6, 16'h6288, 16'h5a68, 16'h6ac9, 16'h5a88, 16'h49e6, 16'h3144, 16'h1881, 16'h3985, 16'h7b6c, 16'h6289, 16'h41c6, 16'h3965, 16'h3124, 16'h3144, 16'h3144, 16'h3164, 16'h3164, 16'h2924, 16'h1061, 16'h820, 16'h820, 16'h1081, 16'h20c2, 16'h293, 16'h3144, 16'h3964, 16'h3985, 16'h41c6, 16'h2924, 16'h41a6, 16'h41c5, 16'h41c5, 16'h41c5, 16'h41c4, 16'h41a4, 16'h41a4, 16'h41a5, 16'h213, 16'h840, 16'h840, 16'h840, 16'h020, 16'h00, 16'h020, 16'h1061, 16'h18a1, 16'h1081, 16'h1061, 16'h1061, 16'h860, 16'h040, 16'h040, 16'h040, 16'h040, 16'h041, 16'h841, 16'h841, 16'h1062, 16'h73b, 16'hde16, 16'hde16, 16'hde16, 16'hde16, 16'hd616, 16'hd616, 16'hd5f6, 16'hd5f6, 16'hd5f6, 16'hd5f5, 16'hd5d5, 16'hd5d5, 16'hd5d5, 16'hd5d5, 16'hcdd5, 16'hcdb5, 16'hcdb5, 16'hcdb5, 16'hcdb5, 16'hcd95, 16'hcd94, 16'hcd94, 16'hcd94, 16'hcd94, 16'hc594, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc573, 16'hc573, 16'hc573, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f2, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacb1, 16'h73b, 16'h2924, 16'h20e2, 16'h20c2, 16'h20c2, 16'h18c2, 16'h1061, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'hb552, 16'hb552, 16'hb552, 16'hb552, 16'hb552, 16'hb552, 16'hb532, 16'had32, 16'had12, 16'had11, 16'had11, 16'hacf1, 16'ha4f1, 16'ha4f1, 16'ha4d1, 16'ha4d0, 16'ha4b0, 16'ha4b0, 16'h9c90, 16'h736b, 16'h20e2, 16'h18a2, 16'h3184, 16'h2123, 16'h1081, 16'h861, 16'h861, 16'h861, 16'h861, 16'h1061, 16'h861, 16'h861, 16'h861, 16'h861, 16'h860, 16'h840, 16'h040, 16'h840, 16'h841, 16'h861, 16'h4a27, 16'h94d, 16'h942e, 16'h942e, 16'h942e, 16'h9c4f, 16'h9c2e, 16'h7b2a, 16'h8bac, 16'h94e, 16'h9c4f, 16'h9c50, 16'h9c4f, 16'h62a9, 16'h20e3, 16'h49e6, 16'h4a7, 16'h6289, 16'h5a68, 16'h4a7, 16'h2923, 16'h1061, 16'h41c6, 16'h7b4b, 16'h5248, 16'h4a6, 16'h49c6, 16'h41c6, 16'h3985, 16'h3164, 16'h3144, 16'h3144, 16'h3144, 16'h20e3, 16'h1081, 16'h840, 16'h840, 16'h840, 16'h841, 16'h1081, 16'h20e3, 16'h213, 16'h2944, 16'h2923, 16'h41c6, 16'h49c5, 16'h41c5, 16'h41c5, 16'h41a4, 16'h41a4, 16'h41a5, 16'h41a4, 16'h293, 16'h841, 16'h840, 16'h840, 16'h020, 16'h00, 16'h820, 16'h1061, 16'h18a1, 16'h1081, 16'h1081, 16'h840, 16'h840, 16'h040, 16'h040, 16'h040, 16'h040, 16'h841, 16'h841, 16'h861, 16'h1062, 16'h73b, 16'hd616, 16'hde16, 16'hd616, 16'hd616, 16'hd5f6, 16'hd5f6, 16'hd5f6, 16'hd5f6, 16'hd5f5, 16'hd5d5, 16'hd5d5, 16'hd5d5, 16'hd5d5, 16'hcdd5, 16'hcdb5, 16'hcdb5, 16'hcdb5, 16'hcdb5, 16'hcdb4, 16'hcd94, 16'hcd94, 16'hcd94, 16'hcd94, 16'hc594, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc573, 16'hc573, 16'hc553, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hac91, 16'h73b, 16'h2923, 16'h20e2, 16'h20c2, 16'h20c2, 16'h20c2, 16'h1061, 16'h020, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'hacf1, 16'hacf1, 16'had11, 16'had11, 16'had32, 16'had32, 16'had12, 16'had32, 16'had11, 16'had11, 16'had11, 16'had11, 16'hacf1, 16'ha4f1, 16'ha4d1, 16'ha4d0, 16'ha4d0, 16'ha4b0, 16'h9cb0, 16'h7b8b, 16'h2123, 16'h18a2, 16'h3185, 16'h213, 16'h1081, 16'h860, 16'h860, 16'h861, 16'h861, 16'h861, 16'h861, 16'h861, 16'h861, 16'h861, 16'h860, 16'h840, 16'h020, 16'h861, 16'h861, 16'h861, 16'h4a27, 16'h94d, 16'h942e, 16'h942e, 16'h942e, 16'h9c4e, 16'h942d, 16'h5247, 16'h732a, 16'h93ed, 16'h94e, 16'h942e, 16'h838c, 16'h49e6, 16'h293, 16'h49e7, 16'h5227, 16'h5a48, 16'h5a68, 16'h49e6, 16'h2923, 16'h18a2, 16'h5248, 16'h73a, 16'h5227, 16'h4a7, 16'h527, 16'h5227, 16'h527, 16'h4a7, 16'h4a7, 16'h49e6, 16'h49e6, 16'h41c6, 16'h41a5, 16'h3164, 16'h20e3, 16'h1081, 16'h840, 16'h840, 16'h840, 16'h861, 16'h1081, 16'h1081, 16'h3984, 16'h39a4, 16'h3984, 16'h41a4, 16'h41a4, 16'h41a5, 16'h39a4, 16'h41a4, 16'h2923, 16'h1081, 16'h1061, 16'h861, 16'h840, 16'h820, 16'h840, 16'h1081, 16'h18a2, 16'h1081, 16'h1081, 16'h1061, 16'h861, 16'h840, 16'h840, 16'h841, 16'h841, 16'h841, 16'h841, 16'h841, 16'h1062, 16'h73b, 16'hd5f6, 16'hd616, 16'hd5f6, 16'hd5f6, 16'hd5f6, 16'hd5f6, 16'hd5f5, 16'hd5f5, 16'hd5d5, 16'hd5d5, 16'hd5d5, 16'hcdd5, 16'hcdd5, 16'hcdb5, 16'hcdb5, 16'hcdb5, 16'hcdb5, 16'hcd94, 16'hcdb4, 16'hcd94, 16'hcd94, 16'hcd94, 16'hc594, 16'hc594, 16'hc574, 16'hc574, 16'hc574, 16'hc573, 16'hc573, 16'hc553, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd32, 16'hbd12, 16'hbd12, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hac90, 16'h73b, 16'h2923, 16'h20e2, 16'h20e2, 16'h20c2, 16'h18c2, 16'h860, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'hacf1, 16'ha4d1, 16'ha4d0, 16'h9cb0, 16'h9c90, 16'h9c90, 16'h9c70, 16'h9c6f, 16'h9c6f, 16'h9c6f, 16'h9c6f, 16'h9c6f, 16'h9c6f, 16'h9c6f, 16'h9c6f, 16'h9c8f, 16'h9c8f, 16'h9c8f, 16'h9c8f, 16'h7b8b, 16'h2923, 16'h18a2, 16'h3184, 16'h213, 16'h1081, 16'h860, 16'h860, 16'h861, 16'h861, 16'h860, 16'h860, 16'h861, 16'h861, 16'h861, 16'h860, 16'h040, 16'h1081, 16'h4a27, 16'h3164, 16'h1061, 16'h4a27, 16'h94d, 16'h942e, 16'h942e, 16'h942d, 16'h9c4e, 16'h942d, 16'h3985, 16'h41a6, 16'h83ad, 16'h94e, 16'h8bed, 16'h73a, 16'h3985, 16'h49e6, 16'h5a68, 16'h5a68, 16'h5a48, 16'h5a48, 16'h41c6, 16'h2924, 16'h293, 16'h5248, 16'h5a68, 16'h527, 16'h4a27, 16'h4a27, 16'h5227, 16'h5227, 16'h5227, 16'h5227, 16'h5227, 16'h49e6, 16'h41c5, 16'h49e6, 16'h4a7, 16'h5227, 16'h41c6, 16'h2924, 16'h18a2, 16'h841, 16'h840, 16'h820, 16'h840, 16'h212, 16'h3123, 16'h3143, 16'h3984, 16'h41a4, 16'h3964, 16'h3143, 16'h3984, 16'h41a4, 16'h3984, 16'h3984, 16'h3164, 16'h3144, 16'h2923, 16'h2923, 16'h2923, 16'h2923, 16'h293, 16'h20e2, 16'h20c2, 16'h18a2, 16'h1081, 16'h1061, 16'h861, 16'h861, 16'h861, 16'h861, 16'h861, 16'h1062, 16'h72eb, 16'hd5f6, 16'hd5f6, 16'hd5f6, 16'hd5f6, 16'hd5f6, 16'hd5f5, 16'hd5f5, 16'hd5d5, 16'hd5d5, 16'hd5d5, 16'hcdd5, 16'hcdb5, 16'hcdb5, 16'hcdb5, 16'hcdb4, 16'hcd94, 16'hcd94, 16'hcd94, 16'hcd94, 16'hcd94, 16'hc594, 16'hc594, 16'hc574, 16'hc574, 16'hc574, 16'hc573, 16'hc573, 16'hc573, 16'hc553, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'ha490, 16'h6aeb, 16'h293, 16'h20e2, 16'h20c2, 16'h20c2, 16'h18c2, 16'h861, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'hbd93, 16'hbd93, 16'hbd73, 16'hb573, 16'hb553, 16'hb553, 16'hb532, 16'had32, 16'had12, 16'hacf1, 16'ha4d1, 16'ha4b0, 16'h9c90, 16'h946f, 16'h944f, 16'h942e, 16'h8ce, 16'h8bed, 16'h8bed, 16'h734a, 16'h2923, 16'h18a2, 16'h3164, 16'h20e2, 16'h861, 16'h861, 16'h860, 16'h861, 16'h860, 16'h860, 16'h860, 16'h860, 16'h860, 16'h860, 16'h860, 16'h040, 16'h1081, 16'h5aa9, 16'h41c5, 16'h1061, 16'h4a7, 16'h94d, 16'h942e, 16'h942e, 16'h942d, 16'h9c4e, 16'h942d, 16'h3984, 16'h18a2, 16'h5228, 16'h8bcd, 16'h8bcd, 16'h527, 16'h41a6, 16'h62a9, 16'h6289, 16'h6289, 16'h5a89, 16'h5248, 16'h4a7, 16'h39a5, 16'h41c6, 16'h5247, 16'h5227, 16'h527, 16'h5227, 16'h5227, 16'h5227, 16'h5227, 16'h5227, 16'h5227, 16'h5227, 16'h41a5, 16'h3164, 16'h3143, 16'h3985, 16'h4a7, 16'h527, 16'h4a6, 16'h41c6, 16'h3144, 16'h3164, 16'h3965, 16'h293, 16'h3123, 16'h41a4, 16'h4184, 16'h3984, 16'h3984, 16'h3984, 16'h3964, 16'h3984, 16'h41a4, 16'h41a4, 16'h41a5, 16'h41c5, 16'h41c5, 16'h41c5, 16'h41c5, 16'h41c5, 16'h41c5, 16'h41c5, 16'h41c5, 16'h41c5, 16'h41a5, 16'h39a5, 16'h3984, 16'h3984, 16'h3164, 16'h3144, 16'h3124, 16'h2923, 16'h2924, 16'h7b4c, 16'hd5f5, 16'hd5f6, 16'hd5f5, 16'hd5f5, 16'hd5f5, 16'hd5d5, 16'hd5d5, 16'hd5d5, 16'hd5d5, 16'hd5b5, 16'hcdb5, 16'hcdb5, 16'hcdb4, 16'hcdb4, 16'hcd94, 16'hcd94, 16'hcd94, 16'hcd94, 16'hcd94, 16'hc594, 16'hc594, 16'hc574, 16'hc574, 16'hc574, 16'hc573, 16'hc573, 16'hc573, 16'hc553, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'ha470, 16'h6aea, 16'h293, 16'h20e2, 16'h20c2, 16'h20c2, 16'h18c2, 16'h841, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'hbd93, 16'hbd93, 16'hbd93, 16'hbd73, 16'hbd73, 16'hb553, 16'hb553, 16'hb552, 16'hb552, 16'hb532, 16'hb532, 16'had32, 16'had12, 16'had12, 16'had11, 16'hacf1, 16'ha4f1, 16'ha4d1, 16'ha4d1, 16'h8cd, 16'h3164, 16'h18a2, 16'h2944, 16'h18e2, 16'h861, 16'h861, 16'h860, 16'h860, 16'h860, 16'h860, 16'h861, 16'h860, 16'h860, 16'h860, 16'h840, 16'h040, 16'h840, 16'h20e3, 16'h18c2, 16'h1061, 16'h4a6, 16'h94d, 16'h94e, 16'h94e, 16'h942e, 16'h9c4e, 16'h942d, 16'h3984, 16'h1041, 16'h20c2, 16'h5a48, 16'h6ac9, 16'h41a5, 16'h5a68, 16'h6aca, 16'h6aaa, 16'h6aaa, 16'h6289, 16'h5228, 16'h41c6, 16'h41a5, 16'h5a48, 16'h5247, 16'h5227, 16'h5227, 16'h5227, 16'h5227, 16'h5227, 16'h5227, 16'h5227, 16'h4a7, 16'h49e6, 16'h41a5, 16'h39a4, 16'h3164, 16'h3985, 16'h49e6, 16'h526, 16'h49e6, 16'h49c5, 16'h527, 16'h73a, 16'h93ed, 16'h7b4b, 16'h6288, 16'h6288, 16'h6288, 16'h6288, 16'h5a68, 16'h5a67, 16'h5a47, 16'h5a47, 16'h5227, 16'h5226, 16'h5226, 16'h4a6, 16'h4a6, 16'h4a6, 16'h49e6, 16'h49e5, 16'h49e5, 16'h49e5, 16'h49e5, 16'h49e5, 16'h49e5, 16'h49e5, 16'h49e6, 16'h49e6, 16'h49e5, 16'h49e5, 16'h49e5, 16'h49e6, 16'h49e6, 16'h8bad, 16'hd5d5, 16'hd5d5, 16'hd5d5, 16'hd5d5, 16'hd5d5, 16'hd5d5, 16'hcdd5, 16'hcdb5, 16'hcdb5, 16'hcdb5, 16'hcdb4, 16'hcdb4, 16'hcd94, 16'hcd94, 16'hcd94, 16'hcd94, 16'hcd94, 16'hc594, 16'hc594, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc573, 16'hc573, 16'hc553, 16'hc553, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'ha470, 16'h6aca, 16'h293, 16'h20e2, 16'h20c2, 16'h20c2, 16'h18a2, 16'h841, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'hbd93, 16'hbd93, 16'hbd73, 16'hbd73, 16'hbd53, 16'hbd53, 16'hb553, 16'hb553, 16'hb553, 16'hb532, 16'hb532, 16'hb532, 16'had32, 16'had12, 16'had12, 16'hacf1, 16'hacf1, 16'hacf1, 16'hacf1, 16'h944e, 16'h3184, 16'h18a2, 16'h2943, 16'h18c2, 16'h861, 16'h861, 16'h840, 16'h860, 16'h860, 16'h860, 16'h860, 16'h840, 16'h840, 16'h860, 16'h860, 16'h840, 16'h840, 16'h861, 16'h861, 16'h1061, 16'h49e6, 16'h94d, 16'h94d, 16'h94e, 16'h942d, 16'h9c4e, 16'h942d, 16'h39a4, 16'h840, 16'h841, 16'h18a2, 16'h3144, 16'h4a7, 16'h6aca, 16'h6aca, 16'h6aea, 16'h6ac9, 16'h5247, 16'h5247, 16'h41c6, 16'h5a48, 16'h6289, 16'h5227, 16'h5227, 16'h5227, 16'h5227, 16'h5227, 16'h5227, 16'h5227, 16'h4a7, 16'h4a7, 16'h41a6, 16'h3985, 16'h3144, 16'h3964, 16'h49e6, 16'h4a6, 16'h51e6, 16'h49c6, 16'h526, 16'h6ac9, 16'h8bac, 16'h8bac, 16'h72e9, 16'h6aa8, 16'h6aa9, 16'h6aa9, 16'h6aa9, 16'h6aa9, 16'h6aa9, 16'h5a68, 16'h5a47, 16'h5a67, 16'h5a67, 16'h5a67, 16'h5a67, 16'h5a68, 16'h6288, 16'h6288, 16'h6288, 16'h6288, 16'h6288, 16'h6288, 16'h5a68, 16'h5a67, 16'h5a67, 16'h5a47, 16'h5247, 16'h5226, 16'h5226, 16'h4a6, 16'h4a6, 16'h527, 16'h8bad, 16'hcdd5, 16'hd5d5, 16'hd5d5, 16'hd5d5, 16'hcdd5, 16'hcdd5, 16'hcdb5, 16'hcdb5, 16'hcdb5, 16'hcdb4, 16'hcdb4, 16'hcd94, 16'hcd94, 16'hcd94, 16'hcd94, 16'hcd94, 16'hc594, 16'hc594, 16'hc594, 16'hc574, 16'hc574, 16'hc574, 16'hc573, 16'hc573, 16'hc573, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f2, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hac90, 16'ha470, 16'h6aca, 16'h293, 16'h20e2, 16'h20c2, 16'h20c2, 16'h18c2, 16'h841, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'hbd73, 16'hbd73, 16'hbd73, 16'hbd53, 16'hbd53, 16'hb553, 16'hb553, 16'hb553, 16'hb553, 16'hb552, 16'hb532, 16'had32, 16'had32, 16'had12, 16'had12, 16'hacf1, 16'hacf1, 16'hacf1, 16'had11, 16'h944e, 16'h3185, 16'h18a2, 16'h213, 16'h10a1, 16'h860, 16'h840, 16'h840, 16'h840, 16'h840, 16'h840, 16'h040, 16'h840, 16'h840, 16'h840, 16'h840, 16'h840, 16'h860, 16'h860, 16'h861, 16'h1061, 16'h49e6, 16'h8bed, 16'h94d, 16'h94d, 16'h94e, 16'h9c4e, 16'h942d, 16'h39a4, 16'h840, 16'h841, 16'h841, 16'h1061, 16'h294, 16'h5a69, 16'h7b6c, 16'h72ea, 16'h5a68, 16'h3965, 16'h5248, 16'h5a48, 16'h62a9, 16'h5248, 16'h5227, 16'h5227, 16'h5227, 16'h5227, 16'h5227, 16'h5227, 16'h5227, 16'h4a7, 16'h41e6, 16'h39a5, 16'h3984, 16'h3164, 16'h41c5, 16'h4a6, 16'h4a6, 16'h49e6, 16'h526, 16'h6aa8, 16'h838b, 16'h838b, 16'h6ac9, 16'h6288, 16'h62a8, 16'h6aa8, 16'h6aa9, 16'h6aa9, 16'h6ac9, 16'h5a67, 16'h527, 16'h526, 16'h526, 16'h526, 16'h4a6, 16'h4a6, 16'h526, 16'h5a47, 16'h5a67, 16'h5a67, 16'h5a47, 16'h5a47, 16'h5a67, 16'h5a67, 16'h5a67, 16'h5a68, 16'h5a88, 16'h5a88, 16'h6288, 16'h62a8, 16'h62a8, 16'h62a8, 16'h6aa9, 16'h94e, 16'hcdd5, 16'hd5d5, 16'hcdd5, 16'hcdd5, 16'hcdb5, 16'hcdb5, 16'hcdb5, 16'hcdb4, 16'hcdb4, 16'hcd94, 16'hcd94, 16'hcd94, 16'hcd94, 16'hc594, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd33, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4d2, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hac90, 16'ha450, 16'h6ac9, 16'h2923, 16'h20e2, 16'h20e2, 16'h20c2, 16'h18a2, 16'h841, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'hbd53, 16'hbd12, 16'hbd52, 16'hbd53, 16'hbd53, 16'hb553, 16'hb553, 16'hb553, 16'hb553, 16'hb553, 16'hb532, 16'hb532, 16'had32, 16'had12, 16'had12, 16'hacf2, 16'hacf1, 16'hacf1, 16'hacf2, 16'h944f, 16'h3985, 16'h18a2, 16'h18e2, 16'h2944, 16'h213, 16'h18c2, 16'h10a1, 16'h1081, 16'h861, 16'h861, 16'h840, 16'h840, 16'h840, 16'h840, 16'h841, 16'h840, 16'h840, 16'h840, 16'h841, 16'h1061, 16'h41c6, 16'h8bed, 16'h94d, 16'h94d, 16'h94d, 16'h9c4e, 16'h942d, 16'h39a4, 16'h840, 16'h841, 16'h841, 16'h841, 16'h1041, 16'h62aa, 16'ha4d0, 16'h6ba, 16'h3165, 16'h20c3, 16'h5a69, 16'h6aea, 16'h6289, 16'h5227, 16'h5227, 16'h5227, 16'h5227, 16'h5227, 16'h5227, 16'h5227, 16'h5227, 16'h4a6, 16'h41c6, 16'h39a5, 16'h3984, 16'h41a5, 16'h49e6, 16'h526, 16'h49e6, 16'h527, 16'h6288, 16'h7b4b, 16'h836b, 16'h62a8, 16'h5a47, 16'h5a47, 16'h5a68, 16'h62a8, 16'h6aa9, 16'h6ac9, 16'h6288, 16'h526, 16'h5227, 16'h5227, 16'h5226, 16'h526, 16'h526, 16'h526, 16'h5227, 16'h5a67, 16'h62a8, 16'h62a8, 16'h5a47, 16'h5a47, 16'h5247, 16'h5227, 16'h5227, 16'h5227, 16'h5227, 16'h5227, 16'h5227, 16'h5227, 16'h5a47, 16'h5a47, 16'h5a48, 16'h8bcd, 16'hcdb5, 16'hcdb5, 16'hcdb5, 16'hcdb5, 16'hcdb5, 16'hcdb4, 16'hcdb4, 16'hcd94, 16'hcd94, 16'hcd94, 16'hcd94, 16'hcd94, 16'hc594, 16'hc594, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc573, 16'hc553, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hacb1, 16'hac90, 16'hac90, 16'ha490, 16'h9c4f, 16'h62a9, 16'h293, 16'h20e2, 16'h20e2, 16'h20c2, 16'h18c2, 16'h841, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'hbd53, 16'hbd12, 16'hbd32, 16'hbd53, 16'hb553, 16'hb553, 16'hb553, 16'hb553, 16'hb552, 16'hb532, 16'hb532, 16'hb532, 16'had12, 16'had12, 16'had12, 16'hacf2, 16'hacf2, 16'hacf2, 16'had11, 16'h946f, 16'h39a5, 16'h18a2, 16'h18c2, 16'h39c5, 16'h39c5, 16'h3185, 16'h2943, 16'h213, 16'h18e3, 16'h18c2, 16'h10a2, 16'h1082, 16'h1081, 16'h1061, 16'h861, 16'h861, 16'h861, 16'h861, 16'h861, 16'h1061, 16'h41a5, 16'h8bed, 16'h94d, 16'h94d, 16'h94d, 16'h9c4e, 16'h942d, 16'h39a5, 16'h840, 16'h840, 16'h841, 16'h841, 16'h1041, 16'h62a9, 16'h8bed, 16'h41c5, 16'h18a2, 16'h18a2, 16'h6aca, 16'h6aea, 16'h5227, 16'h5227, 16'h5227, 16'h5227, 16'h5227, 16'h5227, 16'h5227, 16'h5227, 16'h4a7, 16'h41c5, 16'h41a5, 16'h41c6, 16'h49e6, 16'h5227, 16'h526, 16'h49e6, 16'h5227, 16'h6288, 16'h7b2a, 16'h7b4b, 16'h6288, 16'h41a5, 16'h3143, 16'h3143, 16'h39a5, 16'h4a27, 16'h5a68, 16'h6aa9, 16'h6ac9, 16'h6ac9, 16'h6aa9, 16'h6aa9, 16'h62a8, 16'h62a8, 16'h6288, 16'h6288, 16'h6288, 16'h62a8, 16'h6ac9, 16'h62a8, 16'h6288, 16'h6288, 16'h5a68, 16'h5a47, 16'h5247, 16'h5a47, 16'h5a47, 16'h5247, 16'h5247, 16'h5a47, 16'h5247, 16'h5a47, 16'h5a48, 16'h8bcd, 16'hcdb4, 16'hcdb5, 16'hcdb5, 16'hcdb4, 16'hcdb4, 16'hcd94, 16'hcd94, 16'hcd94, 16'hcd94, 16'hcd94, 16'hcd94, 16'hc594, 16'hc594, 16'hc594, 16'hc574, 16'hc574, 16'hc574, 16'hc573, 16'hc573, 16'hc573, 16'hc553, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hacb0, 16'hacb0, 16'hac90, 16'ha490, 16'ha470, 16'h9c4f, 16'h6289, 16'h28e3, 16'h20e2, 16'h20c2, 16'h20c2, 16'h18a2, 16'h840, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'hbd73, 16'hbd73, 16'hbd53, 16'hbd53, 16'hb553, 16'hb553, 16'hb553, 16'hb553, 16'hb553, 16'hb532, 16'hb532, 16'hb532, 16'had32, 16'had12, 16'had12, 16'had12, 16'hacf1, 16'hacf2, 16'had12, 16'h9c6f, 16'h39a5, 16'h18a2, 16'h18a2, 16'h3185, 16'h39a5, 16'h3184, 16'h2943, 16'h213, 16'h20e3, 16'h18c2, 16'h18a2, 16'h1082, 16'h1081, 16'h1081, 16'h1061, 16'h861, 16'h861, 16'h861, 16'h840, 16'h1061, 16'h41c6, 16'h8bed, 16'h94d, 16'h94d, 16'h94d, 16'h942e, 16'h942d, 16'h41c5, 16'h840, 16'h840, 16'h840, 16'h840, 16'h841, 16'h3985, 16'h4a6, 16'h18a2, 16'h1041, 16'h1061, 16'h5227, 16'h5a88, 16'h4a7, 16'h5227, 16'h5227, 16'h5247, 16'h5247, 16'h5247, 16'h5248, 16'h5248, 16'h5227, 16'h4a7, 16'h5227, 16'h5227, 16'h5227, 16'h5247, 16'h5227, 16'h5a47, 16'h6aa8, 16'h7b4a, 16'h7b4b, 16'h6ac9, 16'h527, 16'h41a5, 16'h3965, 16'h2923, 16'h20e3, 16'h41c6, 16'h5a48, 16'h6288, 16'h6288, 16'h62a8, 16'h62a8, 16'h62a8, 16'h6ac9, 16'h6ac9, 16'h6ae9, 16'h6ae9, 16'h6ae9, 16'h6ae9, 16'h6ac9, 16'h6ac9, 16'h6ac9, 16'h6ae9, 16'h6ac9, 16'h6ac9, 16'h6ac9, 16'h6ac9, 16'h6aa9, 16'h62a8, 16'h62a8, 16'h62a8, 16'h62a8, 16'h6288, 16'h6288, 16'h93ed, 16'hcd94, 16'hcdb4, 16'hcdb4, 16'hcdb4, 16'hcd94, 16'hcd94, 16'hcd94, 16'hcd94, 16'hcd94, 16'hcd94, 16'hc594, 16'hc594, 16'hc574, 16'hc574, 16'hc574, 16'hc573, 16'hc573, 16'hc573, 16'hc553, 16'hc553, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd12, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hb512, 16'hb512, 16'hbd12, 16'hb512, 16'hb4f2, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd0, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'h9c4f, 16'h6289, 16'h293, 16'h20e2, 16'h20c2, 16'h20c2, 16'h18a2, 16'h840, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'hbd73, 16'hbd73, 16'hbd53, 16'hb553, 16'hb553, 16'hb553, 16'hb553, 16'hb553, 16'hb553, 16'hb533, 16'hb532, 16'hb532, 16'had32, 16'had12, 16'had12, 16'had12, 16'hacf2, 16'hacf2, 16'had12, 16'h9c8f, 16'h39a5, 16'h10a2, 16'h18c2, 16'h3184, 16'h39a5, 16'h3164, 16'h2943, 16'h213, 16'h20e3, 16'h18c2, 16'h18a2, 16'h1081, 16'h1081, 16'h1081, 16'h1061, 16'h861, 16'h861, 16'h841, 16'h840, 16'h1061, 16'h41c6, 16'h8bcc, 16'h93ed, 16'h94d, 16'h94d, 16'h942e, 16'h942d, 16'h41c5, 16'h840, 16'h840, 16'h841, 16'h840, 16'h840, 16'h1041, 16'h1061, 16'h840, 16'h840, 16'h820, 16'h1061, 16'h18a2, 16'h18a2, 16'h20e2, 16'h293, 16'h3144, 16'h3964, 16'h3985, 16'h41a5, 16'h49c6, 16'h4a6, 16'h4a27, 16'h5247, 16'h5247, 16'h5a47, 16'h5a47, 16'h5a47, 16'h6ac9, 16'h7b6b, 16'h7b4a, 16'h6ac9, 16'h6aa9, 16'h5a48, 16'h5a48, 16'h5a67, 16'h5a47, 16'h5227, 16'h62a8, 16'h6ac9, 16'h6ac9, 16'h6ac9, 16'h6ac9, 16'h6aa9, 16'h62a8, 16'h62a8, 16'h62a9, 16'h6ae9, 16'h6ae9, 16'h6ae9, 16'h6ae9, 16'h6ae9, 16'h6ae9, 16'h6ae9, 16'h6ae9, 16'h6ae9, 16'h6ae9, 16'h6aea, 16'h6aea, 16'h6ae9, 16'h6ae9, 16'h72e9, 16'h6ae9, 16'h6ae9, 16'h72e9, 16'h72ea, 16'h9c2e, 16'hcd94, 16'hcdb4, 16'hcdb4, 16'hcd94, 16'hcd94, 16'hcd94, 16'hcd94, 16'hcd94, 16'hc594, 16'hc594, 16'hc594, 16'hc574, 16'hc574, 16'hc574, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc553, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb0, 16'hacd0, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'hac90, 16'hac90, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'h9c4f, 16'h6288, 16'h213, 16'h20e2, 16'h20e2, 16'h20c2, 16'h18a2, 16'h840, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'hbd73, 16'hbd73, 16'hbd53, 16'hbd53, 16'hb553, 16'hb553, 16'hb553, 16'hb553, 16'hb553, 16'hb553, 16'hb532, 16'hb532, 16'had32, 16'had12, 16'had12, 16'hacf2, 16'hacf2, 16'hacf2, 16'had12, 16'h9c90, 16'h39a5, 16'h10a1, 16'h18c2, 16'h2964, 16'h3185, 16'h3164, 16'h2923, 16'h213, 16'h20e3, 16'h18c2, 16'h18a2, 16'h1082, 16'h1081, 16'h1081, 16'h1061, 16'h861, 16'h861, 16'h861, 16'h841, 16'h1082, 16'h49e8, 16'h8bcd, 16'h8bed, 16'h93ed, 16'h93ed, 16'h942e, 16'h942d, 16'h41c5, 16'h840, 16'h840, 16'h840, 16'h840, 16'h840, 16'h840, 16'h840, 16'h840, 16'h840, 16'h820, 16'h820, 16'h840, 16'h840, 16'h840, 16'h820, 16'h820, 16'h840, 16'h840, 16'h840, 16'h841, 16'h1041, 16'h1061, 16'h1061, 16'h1882, 16'h1882, 16'h18a2, 16'h49a6, 16'h836b, 16'h7b6b, 16'h6ac9, 16'h6aa9, 16'h6aa9, 16'h6aa9, 16'h6aa9, 16'h6ac9, 16'h6ac9, 16'h6ac9, 16'h6ac9, 16'h6ae9, 16'h6ac9, 16'h6ae9, 16'h6ae9, 16'h6ae9, 16'h6ae9, 16'h6ae9, 16'h6ae9, 16'h6ae9, 16'h6ae9, 16'h6ae9, 16'h6ae9, 16'h6ae9, 16'h6ae9, 16'h6ae9, 16'h6ae9, 16'h6ae9, 16'h6ae9, 16'h6aea, 16'h6aea, 16'h6aea, 16'h6ae9, 16'h72e9, 16'h72e9, 16'h72e9, 16'h72ea, 16'h73a, 16'h9c2e, 16'hc594, 16'hcd94, 16'hcd94, 16'hcd94, 16'hcd94, 16'hcd94, 16'hc594, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc573, 16'hc573, 16'hc553, 16'hc553, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'hac90, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'h9c2e, 16'h5a88, 16'h293, 16'h20e2, 16'h20c2, 16'h18c2, 16'h18a1, 16'h840, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'hbd73, 16'hbd53, 16'hbd53, 16'hbd53, 16'hb553, 16'hb553, 16'hb553, 16'hb553, 16'hb553, 16'hb553, 16'hb532, 16'hb532, 16'had32, 16'had12, 16'had12, 16'hacf2, 16'hacf1, 16'hacf1, 16'had12, 16'h9c90, 16'h39a5, 16'h10a1, 16'h18a2, 16'h2944, 16'h3184, 16'h2944, 16'h2123, 16'h213, 16'h20e3, 16'h18c2, 16'h10a2, 16'h1082, 16'h1081, 16'h1081, 16'h861, 16'h861, 16'h861, 16'h1061, 16'h294, 16'h2969, 16'h5a8c, 16'h8bcd, 16'h8bed, 16'h8bed, 16'h8bed, 16'h942d, 16'h942d, 16'h41c5, 16'h840, 16'h840, 16'h840, 16'h840, 16'h840, 16'h840, 16'h840, 16'h840, 16'h820, 16'h840, 16'h840, 16'h820, 16'h820, 16'h820, 16'h820, 16'h820, 16'h820, 16'h820, 16'h820, 16'h820, 16'h840, 16'h840, 16'h840, 16'h840, 16'h840, 16'h1041, 16'h6288, 16'h838b, 16'h6ac9, 16'h62a8, 16'h6288, 16'h6aa9, 16'h6aa9, 16'h6ac9, 16'h6ac9, 16'h6ac9, 16'h6ac9, 16'h6ac9, 16'h6ac9, 16'h6ae9, 16'h6ae9, 16'h6ae9, 16'h6ae9, 16'h6ae9, 16'h6ae9, 16'h6ae9, 16'h6ae9, 16'h6ae9, 16'h6ae9, 16'h6ae9, 16'h6ae9, 16'h6ae9, 16'h6ae9, 16'h6ae9, 16'h6aea, 16'h6aea, 16'h6aea, 16'h6aea, 16'h72e9, 16'h72e9, 16'h72e9, 16'h72e9, 16'h72e9, 16'h72ea, 16'h73a, 16'h9c2e, 16'hc594, 16'hcd94, 16'hcd94, 16'hc594, 16'hc594, 16'hc594, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc573, 16'hc573, 16'hc573, 16'hc553, 16'hc553, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'hac90, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'h9c2e, 16'h5a68, 16'h213, 16'h20e2, 16'h20c2, 16'h20c2, 16'h18c1, 16'h840, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'hbd73, 16'hbd73, 16'hbd73, 16'hb553, 16'hb553, 16'hb553, 16'hb553, 16'hb553, 16'hb553, 16'hb553, 16'hb532, 16'hb532, 16'had32, 16'had12, 16'had12, 16'hacf2, 16'hacf2, 16'ha4f1, 16'h9cb0, 16'h946f, 16'h39a5, 16'h1081, 16'h10a1, 16'h2944, 16'h3164, 16'h2944, 16'h2123, 16'h213, 16'h18e2, 16'h18c2, 16'h10a2, 16'h1082, 16'h1081, 16'h1061, 16'h861, 16'h861, 16'h861, 16'h214, 16'h5a89, 16'h42c, 16'h5a8d, 16'h83cd, 16'h8bed, 16'h8bed, 16'h8bed, 16'h94e, 16'h942d, 16'h41e5, 16'h840, 16'h840, 16'h840, 16'h841, 16'h840, 16'h840, 16'h820, 16'h820, 16'h820, 16'h820, 16'h820, 16'h840, 16'h820, 16'h820, 16'h820, 16'h820, 16'h820, 16'h820, 16'h820, 16'h820, 16'h820, 16'h820, 16'h840, 16'h840, 16'h840, 16'h1061, 16'h6ac9, 16'h6ae9, 16'h62a9, 16'h6268, 16'h5a47, 16'h62a8, 16'h6aa9, 16'h6ac9, 16'h6ac9, 16'h6ac9, 16'h6ac9, 16'h6ac9, 16'h6ac9, 16'h6ae9, 16'h6ae9, 16'h6ae9, 16'h6ae9, 16'h6ae9, 16'h6ae9, 16'h6ae9, 16'h6ae9, 16'h6ae9, 16'h6ae9, 16'h6ae9, 16'h6ae9, 16'h6ae9, 16'h6ae9, 16'h6ae9, 16'h6ae9, 16'h6aea, 16'h6ae9, 16'h6aea, 16'h72ea, 16'h6ae9, 16'h72e9, 16'h72e9, 16'h72e9, 16'h72ea, 16'h73a, 16'h9c2e, 16'hc594, 16'hcd94, 16'hc594, 16'hc594, 16'hc594, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc553, 16'hc553, 16'hc553, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f2, 16'hb4d2, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'h9c2e, 16'h5a68, 16'h20e3, 16'h20c2, 16'h20c2, 16'h20c1, 16'h18c1, 16'h841, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'hbd73, 16'hbd73, 16'hbd73, 16'hb573, 16'hb553, 16'hb553, 16'hb553, 16'hb553, 16'hb553, 16'hb533, 16'hb512, 16'had12, 16'had32, 16'had12, 16'had12, 16'hacf1, 16'hacf1, 16'h9c90, 16'h5268, 16'h41e6, 16'h213, 16'h1081, 16'h1081, 16'h2923, 16'h3164, 16'h2944, 16'h2123, 16'h20e3, 16'h18e3, 16'h18c2, 16'h10a2, 16'h1082, 16'h1081, 16'h1061, 16'h861, 16'h861, 16'h861, 16'h1082, 16'h2966, 16'h39eb, 16'h524b, 16'h83cd, 16'h8bed, 16'h8bed, 16'h8bed, 16'h94d, 16'h942d, 16'h49e5, 16'h1040, 16'h840, 16'h841, 16'h841, 16'h820, 16'h840, 16'h840, 16'h820, 16'h840, 16'h840, 16'h840, 16'h820, 16'h820, 16'h820, 16'h820, 16'h820, 16'h820, 16'h820, 16'h840, 16'h820, 16'h820, 16'h840, 16'h840, 16'h840, 16'h840, 16'h1061, 16'h5a88, 16'h6ac9, 16'h62a9, 16'h62a9, 16'h5226, 16'h49e5, 16'h49e5, 16'h49e5, 16'h4a6, 16'h5226, 16'h5a67, 16'h5a88, 16'h62a9, 16'h62c9, 16'h6ae9, 16'h6ae9, 16'h6aea, 16'h6aea, 16'h6aea, 16'h6aea, 16'h6ae9, 16'h6ae9, 16'h6ae9, 16'h6ae9, 16'h6ae9, 16'h6aea, 16'h6ae9, 16'h6ae9, 16'h6ae9, 16'h6aea, 16'h6ae9, 16'h6aea, 16'h6aea, 16'h6ae9, 16'h6ae9, 16'h6aea, 16'h6ae9, 16'h72e9, 16'h73a, 16'h942e, 16'hc574, 16'hc594, 16'hc594, 16'hc594, 16'hc594, 16'hc574, 16'hc574, 16'hc574, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc553, 16'hc553, 16'hc553, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hbd12, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha46f, 16'h9ce, 16'h5a48, 16'h20e3, 16'h20c2, 16'h20c2, 16'h20c2, 16'h18a1, 16'h840, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'hbd73, 16'hbd73, 16'hbd73, 16'hb573, 16'hb553, 16'hb553, 16'hb553, 16'hb553, 16'hb533, 16'hb532, 16'hacf2, 16'hacf2, 16'had12, 16'had12, 16'hacf1, 16'hacd1, 16'hacf1, 16'h9c8f, 16'h39a5, 16'h18c2, 16'h18c2, 16'h861, 16'h1061, 16'h213, 16'h2964, 16'h2944, 16'h213, 16'h20e3, 16'h18e2, 16'h18c2, 16'h10a2, 16'h1082, 16'h1081, 16'h1061, 16'h861, 16'h861, 16'h861, 16'h861, 16'h882, 16'h196, 16'h41a8, 16'h83ac, 16'h8bed, 16'h8bed, 16'h8bed, 16'h94e, 16'h94d, 16'h49e5, 16'h841, 16'h840, 16'h840, 16'h841, 16'h840, 16'h840, 16'h840, 16'h840, 16'h820, 16'h820, 16'h820, 16'h820, 16'h820, 16'h820, 16'h820, 16'h820, 16'h820, 16'h820, 16'h820, 16'h820, 16'h820, 16'h840, 16'h820, 16'h821, 16'h1041, 16'h3985, 16'h62a9, 16'h62a9, 16'h62a9, 16'h41c5, 16'h3143, 16'h4183, 16'h3963, 16'h3963, 16'h3943, 16'h3963, 16'h49e5, 16'h4a7, 16'h4a48, 16'h5a89, 16'h62ca, 16'h62ea, 16'h6bb, 16'h732b, 16'h732b, 16'h732b, 16'h6bb, 16'h6ba, 16'h6bb, 16'h6ba, 16'h6aea, 16'h6aea, 16'h6aea, 16'h6ae9, 16'h6aca, 16'h6aca, 16'h6ae9, 16'h6aea, 16'h6aea, 16'h6ae9, 16'h6aea, 16'h6aea, 16'h6ba, 16'h73a, 16'h73a, 16'h94e, 16'hc574, 16'hc594, 16'hc594, 16'hc594, 16'hc594, 16'hc574, 16'hc574, 16'hc574, 16'hc573, 16'hc573, 16'hc573, 16'hc553, 16'hc553, 16'hc553, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hbd12, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f2, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd0, 16'hacb0, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'hac90, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha44f, 16'ha44f, 16'h9ce, 16'h5a48, 16'h20e3, 16'h20c2, 16'h20c2, 16'h20c2, 16'h18a1, 16'h840, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'hbd53, 16'hbd53, 16'hbd73, 16'hb553, 16'hb553, 16'hb553, 16'hb553, 16'hb553, 16'hb533, 16'hb532, 16'had12, 16'had12, 16'hacf2, 16'hacb1, 16'hac91, 16'hac90, 16'hacb1, 16'h9c4f, 16'h41c5, 16'h10a2, 16'h18c2, 16'h1081, 16'h1082, 16'h213, 16'h2944, 16'h2924, 16'h213, 16'h20e3, 16'h18e2, 16'h18c2, 16'h10a2, 16'h1082, 16'h1081, 16'h1061, 16'h1061, 16'h861, 16'h861, 16'h861, 16'h861, 16'h20e3, 16'h527, 16'h83ac, 16'h8bcd, 16'h8bcd, 16'h8bcd, 16'h94d, 16'h94d, 16'h49e5, 16'h840, 16'h840, 16'h840, 16'h840, 16'h840, 16'h840, 16'h840, 16'h841, 16'h840, 16'h820, 16'h820, 16'h820, 16'h820, 16'h820, 16'h840, 16'h840, 16'h820, 16'h820, 16'h820, 16'h820, 16'h820, 16'h820, 16'h821, 16'h1041, 16'h3985, 16'h62a9, 16'h62a9, 16'h62a8, 16'h41a5, 16'h1881, 16'h2922, 16'h4184, 16'h3963, 16'h3963, 16'h3943, 16'h3963, 16'h49e5, 16'h4a7, 16'h5249, 16'h5a89, 16'h62ea, 16'h6bb, 16'h732c, 16'h734d, 16'h734c, 16'h734c, 16'h734c, 16'h732c, 16'h732c, 16'h6b2c, 16'h6bb, 16'h6bb, 16'h6aea, 16'h62ca, 16'h62a9, 16'h6289, 16'h62a9, 16'h62aa, 16'h62ca, 16'h62ca, 16'h6aca, 16'h6aea, 16'h6ba, 16'h6ba, 16'h6bb, 16'h94e, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc573, 16'hc573, 16'hc573, 16'hc553, 16'hc553, 16'hc553, 16'hc553, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hbd12, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f2, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'hac90, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c50, 16'h94e, 16'h5a48, 16'h28e3, 16'h20c2, 16'h20c2, 16'h18c2, 16'h18a1, 16'h840, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'hbd53, 16'hbd32, 16'hbd12, 16'hb532, 16'hb553, 16'hb553, 16'hb553, 16'hb553, 16'hb533, 16'hb533, 16'hb533, 16'had32, 16'hb512, 16'hacb1, 16'hacd2, 16'hacd1, 16'hac90, 16'h9c6f, 16'h41c6, 16'h1081, 16'h1082, 16'h1082, 16'h1082, 16'h213, 16'h2944, 16'h2124, 16'h213, 16'h18e3, 16'h18e2, 16'h18c2, 16'h10a2, 16'h1082, 16'h1081, 16'h1061, 16'h1061, 16'h1061, 16'h861, 16'h841, 16'h861, 16'h213, 16'h6aaa, 16'h8bad, 16'h8bcd, 16'h8bcd, 16'h8bcd, 16'h93ed, 16'h94d, 16'h49e5, 16'h840, 16'h840, 16'h840, 16'h840, 16'h841, 16'h841, 16'h841, 16'h841, 16'h841, 16'h841, 16'h821, 16'h820, 16'h820, 16'h820, 16'h840, 16'h840, 16'h840, 16'h820, 16'h840, 16'h820, 16'h820, 16'h820, 16'h820, 16'h1041, 16'h3124, 16'h3985, 16'h41c6, 16'h3985, 16'h20a2, 16'h1061, 16'h2922, 16'h3984, 16'h3963, 16'h3963, 16'h3963, 16'h3963, 16'h49e6, 16'h4a28, 16'h5269, 16'h5aaa, 16'h6bb, 16'h734c, 16'h736d, 16'h7b6d, 16'h736d, 16'h734d, 16'h734c, 16'h734c, 16'h734c, 16'h732c, 16'h6bb, 16'h6bb, 16'h6aeb, 16'h62ca, 16'h62ca, 16'h62aa, 16'h62aa, 16'h62aa, 16'h62ca, 16'h62cb, 16'h62cb, 16'h62eb, 16'h6bb, 16'h6bb, 16'h6bb, 16'h942f, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc573, 16'hc573, 16'hc573, 16'hc553, 16'hc553, 16'hc553, 16'hc553, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha46f, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h94e, 16'h5248, 16'h20e3, 16'h20c2, 16'h20c2, 16'h18c2, 16'h18a2, 16'h841, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'hbd73, 16'hbd73, 16'hbd33, 16'hbd32, 16'hbd53, 16'hb553, 16'hb512, 16'hb532, 16'hb512, 16'hb512, 16'had32, 16'had32, 16'had12, 16'hacb1, 16'had12, 16'hacd1, 16'hacb1, 16'h9cb0, 16'h41e6, 16'h1082, 16'h1081, 16'h1082, 16'h2082, 16'h314, 16'h2944, 16'h2124, 16'h213, 16'h18e3, 16'h18e2, 16'h18c2, 16'h10a2, 16'h10a2, 16'h1081, 16'h1081, 16'h1061, 16'h1061, 16'h861, 16'h841, 16'h840, 16'h1881, 16'h6ac9, 16'h838c, 16'h83ac, 16'h83ac, 16'h8bcc, 16'h8bed, 16'h94d, 16'h4a6, 16'h18a1, 16'h18a2, 16'h1081, 16'h1061, 16'h1061, 16'h1041, 16'h1041, 16'h841, 16'h841, 16'h841, 16'h841, 16'h840, 16'h821, 16'h820, 16'h840, 16'h840, 16'h820, 16'h840, 16'h820, 16'h820, 16'h841, 16'h840, 16'h841, 16'h821, 16'h821, 16'h841, 16'h1041, 16'h1041, 16'h1041, 16'h1041, 16'h20e2, 16'h3143, 16'h3143, 16'h3143, 16'h3143, 16'h3963, 16'h49e5, 16'h4a28, 16'h5269, 16'h62cb, 16'h734c, 16'h736d, 16'h7b6d, 16'h7b6d, 16'h7b6d, 16'h7b6d, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h6b2b, 16'h6aeb, 16'h6aeb, 16'h6aeb, 16'h6aeb, 16'h62ca, 16'h62ca, 16'h62cb, 16'h62cb, 16'h62eb, 16'h62eb, 16'h62eb, 16'h6bb, 16'h6bb, 16'h6bc, 16'h942f, 16'hc573, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc573, 16'hc573, 16'hc573, 16'hc553, 16'hc553, 16'hc553, 16'hc553, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha44f, 16'ha450, 16'ha450, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h94e, 16'h5247, 16'h20e3, 16'h20e2, 16'h20c2, 16'h18c2, 16'h18a2, 16'h840, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'hb553, 16'hb573, 16'hbd33, 16'hbd13, 16'hbd53, 16'hb553, 16'hb553, 16'hb532, 16'hb512, 16'hb533, 16'had33, 16'had32, 16'hacf2, 16'hac91, 16'hacf2, 16'hacd1, 16'hacb1, 16'ha4b1, 16'h4a6, 16'h10a1, 16'h1081, 16'h1882, 16'h38c3, 16'h3924, 16'h3164, 16'h2944, 16'h213, 16'h18e3, 16'h18e2, 16'h18c2, 16'h10a2, 16'h10a2, 16'h1082, 16'h1081, 16'h1062, 16'h1081, 16'h20e3, 16'h2944, 16'h3164, 16'h525, 16'h8b89, 16'h6aa8, 16'h62a9, 16'h6ac9, 16'h739, 16'h7b4b, 16'h8bcc, 16'h5246, 16'h41c5, 16'h5226, 16'h5226, 16'h5226, 16'h5226, 16'h4a26, 16'h4a6, 16'h49e6, 16'h41c5, 16'h39a5, 16'h3984, 16'h3164, 16'h3144, 16'h293, 16'h20e3, 16'h20c2, 16'h18a2, 16'h1881, 16'h1081, 16'h1061, 16'h1061, 16'h1041, 16'h841, 16'h841, 16'h841, 16'h841, 16'h841, 16'h1041, 16'h1041, 16'h841, 16'h1041, 16'h1881, 16'h1881, 16'h1881, 16'h20a1, 16'h20a2, 16'h293, 16'h41e7, 16'h5a89, 16'h6bb, 16'h7b6d, 16'h7b6d, 16'h7b8d, 16'h7b8d, 16'h7b6d, 16'h7b6d, 16'h736c, 16'h734c, 16'h734c, 16'h734c, 16'h6b2b, 16'h6bb, 16'h6bb, 16'h6bb, 16'h6aeb, 16'h6bb, 16'h6bb, 16'h62eb, 16'h62eb, 16'h6aeb, 16'h62eb, 16'h62eb, 16'h6bb, 16'h6bb, 16'h6bc, 16'h942f, 16'hc573, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc573, 16'hc573, 16'hc553, 16'hc553, 16'hc553, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f2, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha46f, 16'ha44f, 16'ha450, 16'ha450, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h93ee, 16'h5227, 16'h20e3, 16'h20e2, 16'h20c2, 16'h18c2, 16'h18a2, 16'h840, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'hb552, 16'hb553, 16'hbd12, 16'hbcf2, 16'hbd33, 16'hb533, 16'hb553, 16'hb553, 16'hb553, 16'hb553, 16'hb532, 16'had32, 16'had12, 16'hacf2, 16'had12, 16'had12, 16'hacf2, 16'ha4b1, 16'h4a6, 16'h1081, 16'h1061, 16'h2082, 16'h48c3, 16'h394, 16'h3185, 16'h2964, 16'h2123, 16'h18e3, 16'h18e3, 16'h18c2, 16'h10a2, 16'h10a2, 16'h1082, 16'h1081, 16'h1082, 16'h1082, 16'h18a2, 16'h10a2, 16'h1081, 16'h20e2, 16'h4a5, 16'h41c6, 16'h39a7, 16'h39c7, 16'h4a8, 16'h7b4b, 16'h6b9, 16'h3144, 16'h20c2, 16'h20c2, 16'h20e3, 16'h20e3, 16'h213, 16'h2923, 16'h3143, 16'h3164, 16'h3964, 16'h3985, 16'h41a5, 16'h41c5, 16'h41e5, 16'h4a6, 16'h4a6, 16'h526, 16'h5226, 16'h4a6, 16'h5226, 16'h4a26, 16'h4a6, 16'h4a6, 16'h49e6, 16'h41c5, 16'h41a5, 16'h39a5, 16'h3984, 16'h3164, 16'h3144, 16'h20e3, 16'h1061, 16'h1881, 16'h1881, 16'h1861, 16'h20a1, 16'h1881, 16'h20c3, 16'h428, 16'h6aeb, 16'h734c, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h7b6d, 16'h7b6d, 16'h736c, 16'h734c, 16'h734c, 16'h734c, 16'h732c, 16'h732c, 16'h734c, 16'h6b2c, 16'h6bb, 16'h6bb, 16'h6bb, 16'h6aeb, 16'h6aeb, 16'h62eb, 16'h62eb, 16'h62eb, 16'h6bb, 16'h6bb, 16'h6bc, 16'h942f, 16'hc573, 16'hc574, 16'hc574, 16'hc573, 16'hc574, 16'hc573, 16'hc573, 16'hc573, 16'hc553, 16'hc553, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha450, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h93ee, 16'h5227, 16'h20e3, 16'h20e2, 16'h20c2, 16'h18c2, 16'h18a1, 16'h840, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'had12, 16'hb532, 16'hb532, 16'hb4f2, 16'hb512, 16'hb533, 16'hb553, 16'hb553, 16'hb553, 16'hb553, 16'hb553, 16'hb533, 16'had33, 16'had32, 16'had32, 16'hb532, 16'hb513, 16'ha4d1, 16'h4a6, 16'h10a2, 16'h1061, 16'h2082, 16'h48c3, 16'h3924, 16'h41e6, 16'h39c5, 16'h2144, 16'h18e3, 16'h18c2, 16'h10a2, 16'h10a2, 16'h1082, 16'h1061, 16'h861, 16'h861, 16'h861, 16'h1081, 16'h861, 16'h840, 16'h861, 16'h213, 16'h2924, 16'h428, 16'h6bc, 16'h62ca, 16'h7b8c, 16'h41e5, 16'h20c2, 16'h18a2, 16'h18a2, 16'h18a2, 16'h18a2, 16'h18a2, 16'h18a2, 16'h18a2, 16'h18a2, 16'h18a2, 16'h18a2, 16'h18a2, 16'h20c2, 16'h18c2, 16'h20c2, 16'h20c2, 16'h20c2, 16'h20c2, 16'h20c3, 16'h20e3, 16'h20e3, 16'h293, 16'h2924, 16'h3164, 16'h3164, 16'h3985, 16'h39a5, 16'h41c5, 16'h49c6, 16'h49e6, 16'h41c5, 16'h312, 16'h3922, 16'h3942, 16'h3942, 16'h4142, 16'h3942, 16'h3944, 16'h5269, 16'h734c, 16'h7b6d, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h7b6d, 16'h736c, 16'h736c, 16'h736c, 16'h734c, 16'h734c, 16'h736d, 16'h7b6d, 16'h732c, 16'h6b2c, 16'h6bb, 16'h6bb, 16'h6aeb, 16'h6aeb, 16'h6aeb, 16'h62eb, 16'h62eb, 16'h6bb, 16'h6bb, 16'h6b2c, 16'h942f, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc553, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f2, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha44f, 16'ha46f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h93ed, 16'h5227, 16'h20e3, 16'h20c2, 16'h20c2, 16'h20c2, 16'h18a1, 16'h820, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'hacd1, 16'hacd2, 16'hb4f2, 16'hb512, 16'hb512, 16'hb553, 16'hb553, 16'hb553, 16'hb553, 16'hb553, 16'hb553, 16'hb553, 16'hb553, 16'hb533, 16'hb533, 16'hb533, 16'hb533, 16'ha4d1, 16'h4a6, 16'h1082, 16'h1081, 16'h2082, 16'h48c3, 16'h393, 16'h3965, 16'h2923, 16'h20e2, 16'h20e3, 16'h10a2, 16'h861, 16'h861, 16'h861, 16'h861, 16'h860, 16'h841, 16'h841, 16'h1061, 16'h1082, 16'h1082, 16'h18a2, 16'h20e3, 16'h213, 16'h5248, 16'h9c6f, 16'h8bcd, 16'h62a9, 16'h293, 16'h18a2, 16'h18a2, 16'h18a2, 16'h18a2, 16'h18a2, 16'h18a2, 16'h18a2, 16'h18a2, 16'h18a2, 16'h18a2, 16'h18a2, 16'h18a2, 16'h18a2, 16'h20a2, 16'h18c2, 16'h18a2, 16'h18a2, 16'h18a2, 16'h18a2, 16'h18a2, 16'h18a2, 16'h18c2, 16'h20c3, 16'h20e3, 16'h213, 16'h20e3, 16'h213, 16'h213, 16'h294, 16'h3964, 16'h3965, 16'h3964, 16'h3944, 16'h3143, 16'h3143, 16'h3143, 16'h3964, 16'h41a6, 16'h62ca, 16'h734d, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h7b6d, 16'h736d, 16'h734d, 16'h736d, 16'h736d, 16'h7b8d, 16'h7b6d, 16'h7b8d, 16'h732c, 16'h6bc, 16'h6bb, 16'h6bb, 16'h6bb, 16'h6bb, 16'h6bb, 16'h62eb, 16'h6bb, 16'h6bc, 16'h6b2b, 16'h732c, 16'h942f, 16'hc573, 16'hc573, 16'hc573, 16'hc574, 16'hc574, 16'hc573, 16'hc573, 16'hc553, 16'hc553, 16'hc553, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha450, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h93ed, 16'h5226, 16'h20e3, 16'h20c2, 16'h20c2, 16'h20c2, 16'h18a1, 16'h840, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'ha4b0, 16'ha4b1, 16'hac91, 16'hb4b1, 16'hb4d2, 16'hb512, 16'hb533, 16'hb553, 16'hb553, 16'hb553, 16'hb553, 16'hb553, 16'hb553, 16'hb553, 16'hb553, 16'hb553, 16'hb553, 16'hacf2, 16'h4a7, 16'h1081, 16'h1081, 16'h2082, 16'h40c3, 16'h3061, 16'h2861, 16'h2061, 16'h2061, 16'h28e3, 16'h20e3, 16'h10a2, 16'h861, 16'h18e3, 16'h18c2, 16'h860, 16'h20e3, 16'h3165, 16'h41c6, 16'h3185, 16'h2944, 16'h20e3, 16'h10a2, 16'h10a2, 16'h41c6, 16'h942e, 16'h62c9, 16'h3144, 16'h18a2, 16'h1881, 16'h1081, 16'h1081, 16'h1082, 16'h1882, 16'h1082, 16'h18a2, 16'h18a2, 16'h18a2, 16'h18a2, 16'h18a2, 16'h1882, 16'h18a2, 16'h20a2, 16'h20c2, 16'h18c2, 16'h18a2, 16'h18a2, 16'h18a2, 16'h18a2, 16'h18a2, 16'h18c2, 16'h20c3, 16'h20e3, 16'h20e3, 16'h20e3, 16'h213, 16'h2924, 16'h41a5, 16'h4a6, 16'h4a6, 16'h49e6, 16'h49e5, 16'h49c6, 16'h49c5, 16'h49e6, 16'h5a27, 16'h5a89, 16'h6b2c, 16'h736d, 16'h7b8d, 16'h7bad, 16'h7bad, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h736d, 16'h736d, 16'h7b6d, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h6b2c, 16'h6b2c, 16'h6b2b, 16'h6b2c, 16'h6bc, 16'h6bb, 16'h6aeb, 16'h62eb, 16'h6bb, 16'h6b2c, 16'h6b2b, 16'h732c, 16'h942f, 16'hc573, 16'hc574, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc553, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha450, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h93ed, 16'h4a6, 16'h20e3, 16'h20c2, 16'h20c2, 16'h20c2, 16'h18a1, 16'h820, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h9c70, 16'h9c90, 16'ha4b1, 16'hacd2, 16'hacf2, 16'had12, 16'hb532, 16'hb533, 16'hb553, 16'hb553, 16'hb553, 16'hb554, 16'hbd74, 16'hbd74, 16'hbd54, 16'hbd54, 16'hb553, 16'had12, 16'h4a27, 16'h1082, 16'h1081, 16'h2082, 16'h40a2, 16'h3061, 16'h2841, 16'h2040, 16'h2061, 16'h28c2, 16'h2944, 16'h18a2, 16'h840, 16'h10a2, 16'h10a2, 16'h861, 16'h5247, 16'h732a, 16'h732a, 16'h6ba, 16'h732a, 16'h41c5, 16'h840, 16'h840, 16'h41c6, 16'h942e, 16'h49e6, 16'h18a2, 16'h1082, 16'h1081, 16'h1061, 16'h1061, 16'h1061, 16'h1061, 16'h1061, 16'h1061, 16'h1081, 16'h1082, 16'h1082, 16'h1882, 16'h1882, 16'h18a2, 16'h18a2, 16'h18a2, 16'h18a2, 16'h18a2, 16'h18a2, 16'h18a2, 16'h18a2, 16'h18a2, 16'h18c2, 16'h18c3, 16'h20e3, 16'h20e3, 16'h20e3, 16'h3124, 16'h41a5, 16'h4a6, 16'h4a6, 16'h4a6, 16'h49e6, 16'h49e6, 16'h49e5, 16'h5227, 16'h5a68, 16'h5a89, 16'h62cb, 16'h734c, 16'h7b6d, 16'h7b8d, 16'h7bad, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h7b6d, 16'h7b6d, 16'h7b6d, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h6b2c, 16'h6b2c, 16'h6b2b, 16'h6b2c, 16'h6b2c, 16'h6bc, 16'h6aeb, 16'h6aeb, 16'h6bb, 16'h732c, 16'h732b, 16'h732c, 16'h942f, 16'hc573, 16'hc574, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc553, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h93cd, 16'h4a6, 16'h20e3, 16'h20c2, 16'h20c2, 16'h18c2, 16'h18a2, 16'h820, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h944f, 16'h9c70, 16'ha4b1, 16'ha4d1, 16'hacf2, 16'had12, 16'hb533, 16'hb533, 16'hb553, 16'hb553, 16'hb533, 16'hbd53, 16'hbd54, 16'hbd74, 16'hbd74, 16'hbd74, 16'hbd74, 16'hb532, 16'h4a27, 16'h1082, 16'h1081, 16'h2082, 16'h40a2, 16'h3061, 16'h2841, 16'h2840, 16'h2040, 16'h2081, 16'h28e2, 16'h1881, 16'h1061, 16'h1061, 16'h841, 16'h1082, 16'h5248, 16'h732a, 16'h732a, 16'h732a, 16'h838b, 16'h4a6, 16'h840, 16'h820, 16'h2944, 16'h5a88, 16'h20e2, 16'h1061, 16'h1061, 16'h1061, 16'h1081, 16'h1061, 16'h1081, 16'h1081, 16'h1082, 16'h1082, 16'h1082, 16'h1082, 16'h1082, 16'h1082, 16'h1882, 16'h18a2, 16'h18a2, 16'h18a2, 16'h18a2, 16'h18a2, 16'h18a2, 16'h18a2, 16'h1882, 16'h18a2, 16'h18a2, 16'h18c2, 16'h20e3, 16'h20e3, 16'h3144, 16'h41c5, 16'h4a6, 16'h4a6, 16'h4a6, 16'h49e6, 16'h49e6, 16'h49e6, 16'h5227, 16'h5268, 16'h5269, 16'h5aaa, 16'h6bc, 16'h736d, 16'h7b8e, 16'h7b8d, 16'h7bad, 16'h7bad, 16'h7b8d, 16'h7b8d, 16'h7b6d, 16'h7b6d, 16'h7b6d, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h6b2c, 16'h6b2c, 16'h6b2c, 16'h6b2c, 16'h6b2c, 16'h6b2c, 16'h6bc, 16'h6bb, 16'h6bb, 16'h732c, 16'h732b, 16'h732b, 16'h942f, 16'hc573, 16'hc574, 16'hc574, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc553, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd52, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha44f, 16'ha450, 16'ha450, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h93cd, 16'h4a6, 16'h20e2, 16'h20e2, 16'h20c2, 16'h20c2, 16'h18a2, 16'h820, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h94f, 16'h9450, 16'h9c90, 16'h9cb1, 16'ha4d1, 16'hacf2, 16'had12, 16'hb533, 16'hb533, 16'hb553, 16'hb513, 16'hbd54, 16'hbd74, 16'hbd74, 16'hbd74, 16'hbd74, 16'hbd94, 16'hb553, 16'h4a27, 16'h1082, 16'h1082, 16'h2082, 16'h40a2, 16'h2861, 16'h2841, 16'h2841, 16'h2040, 16'h2040, 16'h2041, 16'h2041, 16'h2061, 16'h2862, 16'h2861, 16'h2882, 16'h5a48, 16'h732a, 16'h732a, 16'h732a, 16'h838b, 16'h4a6, 16'h840, 16'h020, 16'h820, 16'h861, 16'h020, 16'h020, 16'h020, 16'h020, 16'h820, 16'h820, 16'h820, 16'h820, 16'h820, 16'h840, 16'h841, 16'h841, 16'h841, 16'h841, 16'h1061, 16'h1061, 16'h1061, 16'h1081, 16'h1081, 16'h1081, 16'h1881, 16'h1881, 16'h1882, 16'h18a2, 16'h18a2, 16'h20c2, 16'h20e3, 16'h3144, 16'h41e6, 16'h526, 16'h4a6, 16'h4a6, 16'h49e6, 16'h49e5, 16'h49e6, 16'h5227, 16'h5268, 16'h5269, 16'h5aaa, 16'h62eb, 16'h6b2c, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h7b6d, 16'h736d, 16'h7b6d, 16'h7b8d, 16'h7b8d, 16'h7bad, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h6b2c, 16'h6b2c, 16'h6b2c, 16'h732c, 16'h6b2c, 16'h6b2b, 16'h6b2b, 16'h6b2b, 16'h6bb, 16'h732c, 16'h732c, 16'h732c, 16'h9c2f, 16'hc573, 16'hc574, 16'hc574, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd52, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hbd12, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha470, 16'ha46f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h93cd, 16'h49e6, 16'h20e2, 16'h20e2, 16'h20c2, 16'h20c2, 16'h18a1, 16'h820, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h8bee, 16'h942f, 16'h9c70, 16'h9c91, 16'ha4d1, 16'hacf2, 16'had12, 16'hb533, 16'hb533, 16'hb553, 16'hbd54, 16'hbd54, 16'hbd54, 16'hc595, 16'hc595, 16'hbd94, 16'hbd94, 16'hb553, 16'h4a27, 16'h1082, 16'h1062, 16'h2082, 16'h40a2, 16'h2861, 16'h2841, 16'h2041, 16'h2040, 16'h2040, 16'h2040, 16'h2020, 16'h2841, 16'h3041, 16'h3061, 16'h30a4, 16'h6269, 16'h732a, 16'h732a, 16'h732a, 16'h838b, 16'h4a26, 16'h840, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h820, 16'h820, 16'h1061, 16'h18a1, 16'h20c1, 16'h20e1, 16'h20e2, 16'h3144, 16'h41c6, 16'h4a27, 16'h5268, 16'h5268, 16'h5268, 16'h5268, 16'h5248, 16'h5228, 16'h5248, 16'h5269, 16'h5269, 16'h5a89, 16'h62ca, 16'h6bb, 16'h734c, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h736d, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h734c, 16'h6b2c, 16'h6b2c, 16'h732c, 16'h6b2c, 16'h6b2b, 16'h6b2b, 16'h6b2b, 16'h6b2c, 16'h732c, 16'h732b, 16'h734c, 16'h9c2f, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc553, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha450, 16'ha44f, 16'ha44f, 16'h9c4f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h93cd, 16'h49e6, 16'h20e2, 16'h20c2, 16'h20c2, 16'h20c2, 16'h18a1, 16'h820, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h8bef, 16'h9430, 16'h9c70, 16'h9c91, 16'ha4d1, 16'ha4f2, 16'had12, 16'hb513, 16'hb533, 16'hb554, 16'hbd54, 16'hbd54, 16'hbd54, 16'hbd74, 16'hbd95, 16'hbd94, 16'hbd94, 16'hb553, 16'h5a69, 16'h20e3, 16'h18a2, 16'h2082, 16'h40a2, 16'h3061, 16'h2841, 16'h2041, 16'h2040, 16'h2040, 16'h2040, 16'h2040, 16'h2841, 16'h3041, 16'h414, 16'h3969, 16'h62cd, 16'h732a, 16'h732a, 16'h732a, 16'h838b, 16'h4a26, 16'h840, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h820, 16'h1060, 16'h18a1, 16'h20c1, 16'h20e2, 16'h20e2, 16'h3164, 16'h4a27, 16'h5269, 16'h5289, 16'h5a89, 16'h5a89, 16'h5a89, 16'h5a89, 16'h5a89, 16'h5a89, 16'h5289, 16'h5289, 16'h5aaa, 16'h62eb, 16'h6b2c, 16'h734d, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h7b6d, 16'h736d, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h7b6d, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h734c, 16'h6b2c, 16'h6b2c, 16'h6b2c, 16'h6b2c, 16'h6b2b, 16'h6b2b, 16'h6b2c, 16'h6b2c, 16'h732c, 16'h732c, 16'h734c, 16'h9c4f, 16'hc573, 16'hc574, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd12, 16'hbd12, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb0, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha48f, 16'ha46f, 16'ha470, 16'ha470, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h8bcd, 16'h49e6, 16'h20e2, 16'h20c2, 16'h20c2, 16'h20c2, 16'h18a1, 16'h820, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h94f, 16'h9450, 16'h9c70, 16'h9cb1, 16'ha4d2, 16'hacf2, 16'hacf2, 16'hb4f2, 16'hb533, 16'hb554, 16'hbd74, 16'hbd74, 16'hbd74, 16'hbd74, 16'hbd95, 16'hbd94, 16'hbd94, 16'hbd94, 16'ha4d2, 16'h9c91, 16'h83ad, 16'h49c6, 16'h413, 16'h3061, 16'h2861, 16'h2841, 16'h2040, 16'h2040, 16'h2041, 16'h2841, 16'h2841, 16'h3062, 16'h4986, 16'h4a2c, 16'h6acc, 16'h732a, 16'h732a, 16'h732a, 16'h838b, 16'h4a26, 16'h840, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h820, 16'h1060, 16'h18a1, 16'h20e2, 16'h20e2, 16'h20e2, 16'h3964, 16'h4a27, 16'h5a89, 16'h5a89, 16'h5aa9, 16'h5aa9, 16'h5aa9, 16'h5aa9, 16'h5aa9, 16'h5aa9, 16'h5aaa, 16'h5aaa, 16'h62ca, 16'h6bb, 16'h6b2c, 16'h7b6d, 16'h7b8d, 16'h7bad, 16'h7b8d, 16'h7b6d, 16'h7b6d, 16'h7b6d, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h7b8e, 16'h7bad, 16'h7b8d, 16'h7b8d, 16'h734c, 16'h732c, 16'h734c, 16'h6b2c, 16'h6b2c, 16'h6b2c, 16'h6b2c, 16'h6b2c, 16'h6b2b, 16'h732c, 16'h732c, 16'h732c, 16'h9c2f, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd12, 16'hbd12, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb0, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha470, 16'ha470, 16'ha44f, 16'ha44f, 16'ha450, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h8bad, 16'h49e6, 16'h20e2, 16'h20c2, 16'h20c2, 16'h18c2, 16'h18a1, 16'h820, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h942f, 16'h9c50, 16'h9c91, 16'ha4b1, 16'ha4d2, 16'hacd2, 16'hacf2, 16'hb513, 16'hb533, 16'hb554, 16'hbd54, 16'hbd74, 16'hbd74, 16'hbd74, 16'hbd94, 16'hbd94, 16'hbd94, 16'hbd94, 16'hc594, 16'hc5b5, 16'hacf1, 16'h5248, 16'h49a5, 16'h40e4, 16'h3062, 16'h2861, 16'h2841, 16'h2841, 16'h2841, 16'h2841, 16'h2841, 16'h2841, 16'h30c4, 16'h3967, 16'h5a69, 16'h732a, 16'h732a, 16'h7b4a, 16'h83ac, 16'h5247, 16'h861, 16'h820, 16'h820, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h820, 16'h820, 16'h820, 16'h1081, 16'h18a1, 16'h20e2, 16'h28e2, 16'h28e2, 16'h3984, 16'h5248, 16'h5a89, 16'h5a89, 16'h5aa9, 16'h5ac9, 16'h5aa9, 16'h5aaa, 16'h5aa9, 16'h5aa9, 16'h5aaa, 16'h62cb, 16'h62eb, 16'h6bc, 16'h734c, 16'h7b8d, 16'h7bad, 16'h7bae, 16'h7bad, 16'h7b8d, 16'h7b6d, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h7bae, 16'h7bae, 16'h7bad, 16'h7b8d, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h732c, 16'h732c, 16'h6b2c, 16'h6b2c, 16'h6b2b, 16'h6b2c, 16'h732c, 16'h734c, 16'h9c4f, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc553, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hacd1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h8bad, 16'h49e6, 16'h20e2, 16'h20c2, 16'h20c2, 16'h18c2, 16'h18a1, 16'h820, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h9c50, 16'h9c91, 16'ha471, 16'ha491, 16'hacd2, 16'hacf2, 16'hb513, 16'hb533, 16'hb533, 16'hb533, 16'hb554, 16'hbd54, 16'hbd74, 16'hbd74, 16'hbd74, 16'hbd74, 16'hbd94, 16'hbd94, 16'hbd94, 16'hc5b5, 16'hacf1, 16'h5248, 16'h5248, 16'h72ea, 16'h6228, 16'h4945, 16'h38c3, 16'h3082, 16'h3062, 16'h2861, 16'h2841, 16'h30a3, 16'h30c3, 16'h38e3, 16'h5a27, 16'h6288, 16'h6ac9, 16'h6ae9, 16'h838b, 16'h5a87, 16'h2923, 16'h3144, 16'h3144, 16'h2944, 16'h2923, 16'h2923, 16'h213, 16'h20e3, 16'h20c2, 16'h18c2, 16'h18a2, 16'h18a2, 16'h1081, 16'h1081, 16'h1061, 16'h1061, 16'h861, 16'h841, 16'h841, 16'h840, 16'h820, 16'h820, 16'h820, 16'h820, 16'h1061, 16'h18a1, 16'h20e2, 16'h292, 16'h292, 16'h3984, 16'h5248, 16'h5a89, 16'h5aa9, 16'h5aaa, 16'h62ca, 16'h62ca, 16'h62ca, 16'h5aaa, 16'h5aaa, 16'h62ca, 16'h62eb, 16'h62eb, 16'h6bb, 16'h734c, 16'h7b8d, 16'h7bae, 16'h7bad, 16'h7bad, 16'h7b6d, 16'h7b6d, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h7bad, 16'h7bae, 16'h7bae, 16'h7bad, 16'h7b8d, 16'h736c, 16'h734c, 16'h734c, 16'h734c, 16'h732c, 16'h6b2c, 16'h6b2c, 16'h6b2b, 16'h6b2b, 16'h734c, 16'h734c, 16'h734b, 16'h9c4f, 16'hc573, 16'hc574, 16'hc574, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc553, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha46f, 16'ha450, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h8bad, 16'h49e5, 16'h20e2, 16'h20c2, 16'h20c2, 16'h18c2, 16'h18a1, 16'h820, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'ha491, 16'ha4b1, 16'hac71, 16'hac92, 16'had13, 16'hb513, 16'hb533, 16'hb534, 16'hb533, 16'hb534, 16'hb554, 16'hb554, 16'hbd54, 16'hbd54, 16'hbd74, 16'hbd74, 16'hbd74, 16'hbd74, 16'hbd74, 16'hbd94, 16'ha4d1, 16'h5268, 16'h5248, 16'h83cd, 16'h9c70, 16'h9c50, 16'h93ee, 16'h836c, 16'h72ca, 16'h51a6, 16'h393, 16'h394, 16'h38e3, 16'h4123, 16'h4984, 16'h4164, 16'h4985, 16'h526, 16'h62a8, 16'h3984, 16'h18a1, 16'h18a2, 16'h18a2, 16'h18a2, 16'h18a2, 16'h18c2, 16'h18c2, 16'h20e2, 16'h213, 16'h293, 16'h293, 16'h2923, 16'h2923, 16'h2943, 16'h2943, 16'h2944, 16'h2944, 16'h2943, 16'h2943, 16'h3143, 16'h2943, 16'h2923, 16'h2923, 16'h213, 16'h18c1, 16'h20c1, 16'h20e2, 16'h292, 16'h292, 16'h3984, 16'h5268, 16'h5aa9, 16'h5aa9, 16'h62ca, 16'h62ca, 16'h62ca, 16'h62ca, 16'h62ca, 16'h62ca, 16'h62eb, 16'h62eb, 16'h62eb, 16'h6b2c, 16'h736d, 16'h7b8d, 16'h7bae, 16'h7bad, 16'h7b8e, 16'h7b6d, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h7bad, 16'h83ae, 16'h83ae, 16'h83ae, 16'h7bad, 16'h7bad, 16'h7b8d, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h6b2c, 16'h6b2c, 16'h6b2c, 16'h6b2b, 16'h6b2b, 16'h732c, 16'h734c, 16'h734c, 16'h9c4f, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc553, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4e, 16'h9c2e, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h8bac, 16'h41c5, 16'h20e2, 16'h20c2, 16'h18c2, 16'h18c2, 16'h18a1, 16'h820, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'hac71, 16'hacd2, 16'hacb2, 16'hb4b2, 16'hb513, 16'hb533, 16'hb534, 16'hb534, 16'hb533, 16'hb534, 16'hb554, 16'hb554, 16'hb554, 16'hb554, 16'hb554, 16'hb554, 16'hb554, 16'hb554, 16'hbd74, 16'hbd74, 16'ha4d1, 16'h5248, 16'h5248, 16'h83ad, 16'h9c90, 16'h9c91, 16'h83ad, 16'h944f, 16'h734b, 16'h4a6, 16'h3124, 16'h3124, 16'h5a47, 16'h6287, 16'h5a26, 16'h4184, 16'h525, 16'h49c4, 16'h49a4, 16'h3963, 16'h3142, 16'h3122, 16'h3122, 16'h292, 16'h292, 16'h292, 16'h20e2, 16'h28e2, 16'h20e2, 16'h20e1, 16'h20c1, 16'h20c2, 16'h20c2, 16'h20c2, 16'h20c2, 16'h20a2, 16'h18a2, 16'h18a1, 16'h18a1, 16'h20c2, 16'h20a2, 16'h18a2, 16'h18a1, 16'h20c2, 16'h20e2, 16'h20e2, 16'h18c2, 16'h18a1, 16'h18a1, 16'h2923, 16'h5268, 16'h5aaa, 16'h5aca, 16'h62ca, 16'h62ea, 16'h62ca, 16'h62ea, 16'h62eb, 16'h62ca, 16'h62ea, 16'h62eb, 16'h6bb, 16'h732c, 16'h7b6d, 16'h7b8d, 16'h7b8e, 16'h7bad, 16'h7bad, 16'h7b6d, 16'h7b6d, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h7bae, 16'h83ae, 16'h83ce, 16'h83ce, 16'h83ae, 16'h7bad, 16'h7b8d, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h732c, 16'h6b2c, 16'h6b2b, 16'h6bb, 16'h6b2c, 16'h734c, 16'h734c, 16'h7b4c, 16'h9c4f, 16'hc573, 16'hc573, 16'hc574, 16'hc574, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc553, 16'hc553, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha46f, 16'ha470, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h8bad, 16'h41c5, 16'h20e2, 16'h20c2, 16'h20c2, 16'h18c2, 16'h18a1, 16'h820, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'hac71, 16'hb4d2, 16'hb4d2, 16'hb4d3, 16'hb513, 16'hb514, 16'hb534, 16'hb534, 16'hb513, 16'hb513, 16'hb534, 16'hb534, 16'hb534, 16'hb533, 16'hb533, 16'hb533, 16'hb533, 16'hb533, 16'hb553, 16'hbd74, 16'ha4d1, 16'h5268, 16'h5248, 16'h7bad, 16'h9c90, 16'h9450, 16'h41e7, 16'h5268, 16'h294, 16'h1881, 16'h1881, 16'h20e3, 16'h6288, 16'h72e9, 16'h5a46, 16'h28e2, 16'h6aea, 16'h41c5, 16'h20a2, 16'h20a1, 16'h18a1, 16'h20a1, 16'h18a2, 16'h18c1, 16'h18c1, 16'h20c2, 16'h3123, 16'h3983, 16'h292, 16'h292, 16'h292, 16'h292, 16'h292, 16'h3122, 16'h3122, 16'h3123, 16'h3122, 16'h3122, 16'h3122, 16'h3122, 16'h3122, 16'h3142, 16'h3942, 16'h3943, 16'h3963, 16'h2923, 16'h20e2, 16'h18c2, 16'h861, 16'h18a2, 16'h4a48, 16'h62ca, 16'h62ca, 16'h62ea, 16'h62ea, 16'h62ea, 16'h62ea, 16'h62ea, 16'h62ca, 16'h62ea, 16'h6bb, 16'h6bb, 16'h734c, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h7bad, 16'h7bad, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h7b8e, 16'h7bae, 16'h7bae, 16'h7bad, 16'h83ce, 16'h83ce, 16'h83ce, 16'h83ad, 16'h7b8d, 16'h7b8d, 16'h734c, 16'h6b2c, 16'h732c, 16'h734c, 16'h6b2b, 16'h6b2c, 16'h6b2b, 16'h6bb, 16'h6bb, 16'h734c, 16'h734c, 16'h734c, 16'h9c4f, 16'hc573, 16'hc574, 16'hc574, 16'hc574, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha470, 16'ha46f, 16'ha46f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h8bad, 16'h41a5, 16'h20e2, 16'h20c2, 16'h20c2, 16'h20c1, 16'h18a1, 16'h820, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'hb4b2, 16'hb4f3, 16'hb4d3, 16'hb4f3, 16'hb513, 16'hb514, 16'hb534, 16'hb534, 16'hb534, 16'hb513, 16'hb533, 16'hb534, 16'hb533, 16'hb533, 16'hb513, 16'hb513, 16'hb533, 16'hb533, 16'hb553, 16'hbd74, 16'ha4d1, 16'h5248, 16'h4a48, 16'h7b8d, 16'h9c70, 16'h62ca, 16'h5269, 16'h7b8d, 16'h5a8a, 16'h4a8, 16'h5a48, 16'h5a67, 16'h7b29, 16'h7b9, 16'h5a47, 16'h20a2, 16'h3985, 16'h18c2, 16'h18c2, 16'h18a2, 16'h18a1, 16'h1081, 16'h1082, 16'h1081, 16'h1081, 16'h1081, 16'h292, 16'h3963, 16'h1881, 16'h1040, 16'h840, 16'h840, 16'h841, 16'h1061, 16'h1061, 16'h1061, 16'h1061, 16'h1061, 16'h1061, 16'h1881, 16'h18a1, 16'h28e1, 16'h4183, 16'h49c4, 16'h3963, 16'h1081, 16'h1081, 16'h1061, 16'h841, 16'h213, 16'h5a89, 16'h6aeb, 16'h6aeb, 16'h6bb, 16'h6bb, 16'h6bb, 16'h6aeb, 16'h62ea, 16'h62ea, 16'h62eb, 16'h6bb, 16'h6b2b, 16'h734c, 16'h7b8d, 16'h7b8d, 16'h7bad, 16'h83ae, 16'h7bad, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h7bae, 16'h7bae, 16'h7bae, 16'h83ae, 16'h83ce, 16'h83ce, 16'h83ce, 16'h83ad, 16'h7b8d, 16'h7b8d, 16'h732c, 16'h6b2c, 16'h732c, 16'h732b, 16'h6b2b, 16'h6b2b, 16'h6b2b, 16'h6bb, 16'h6b2b, 16'h734c, 16'h734c, 16'h734c, 16'h9c2f, 16'hc573, 16'hc594, 16'hc574, 16'hc574, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc553, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb0, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha46f, 16'ha470, 16'ha46f, 16'ha470, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h8bac, 16'h41a5, 16'h20e2, 16'h20c2, 16'h20c2, 16'h20c2, 16'h18a1, 16'h820, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'hb4b2, 16'hb4f3, 16'hb4f3, 16'hbcf3, 16'hbd13, 16'hb534, 16'hb533, 16'hb513, 16'hb513, 16'hacf3, 16'hacf2, 16'hb513, 16'hb513, 16'had13, 16'had13, 16'had13, 16'had13, 16'hb513, 16'hb533, 16'hb554, 16'ha4b1, 16'h5248, 16'h4a27, 16'h6b2b, 16'h62ca, 16'h41c6, 16'h7b8d, 16'h942f, 16'h9c70, 16'h8bce, 16'h73a, 16'h6ac9, 16'h834a, 16'h72e9, 16'h5a47, 16'h20a1, 16'h1061, 16'h1061, 16'h18c2, 16'h213, 16'h2924, 16'h213, 16'h20e3, 16'h213, 16'h213, 16'h20e2, 16'h3143, 16'h4183, 16'h1881, 16'h1060, 16'h1060, 16'h1060, 16'h1060, 16'h1060, 16'h1061, 16'h1061, 16'h1060, 16'h1060, 16'h1060, 16'h1881, 16'h20c1, 16'h20c1, 16'h4184, 16'h49c4, 16'h3963, 16'h840, 16'h020, 16'h020, 16'h841, 16'h2945, 16'h5aa9, 16'h6bb, 16'h6bb, 16'h6bb, 16'h6b2b, 16'h6bb, 16'h6bb, 16'h6aeb, 16'h62eb, 16'h6bb, 16'h6bb, 16'h6b2c, 16'h736c, 16'h7bad, 16'h7bad, 16'h83ad, 16'h83ae, 16'h7bae, 16'h7b8d, 16'h7b8d, 16'h7bad, 16'h83ae, 16'h7bae, 16'h7bae, 16'h83ae, 16'h83ce, 16'h83ce, 16'h83cd, 16'h7bad, 16'h7bad, 16'h7b8d, 16'h734c, 16'h6b2b, 16'h6b2c, 16'h6b2c, 16'h6b2b, 16'h6bb, 16'h6bb, 16'h6bb, 16'h6bb, 16'h732c, 16'h734c, 16'h734d, 16'h9c4f, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc553, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb0, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha46f, 16'ha470, 16'ha470, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h8bac, 16'h41a5, 16'h20e2, 16'h20c2, 16'h20c2, 16'h20c2, 16'h18a1, 16'h820, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'hb4f3, 16'hbcf3, 16'hbd14, 16'hbcf3, 16'hb4f3, 16'hb534, 16'hb533, 16'had13, 16'hacf3, 16'hacf3, 16'hacd3, 16'hacf3, 16'hacf3, 16'hacf3, 16'hacf3, 16'hacf3, 16'hacf3, 16'hacd2, 16'ha4d2, 16'ha4b1, 16'h838c, 16'h41c6, 16'h3985, 16'h3985, 16'h3145, 16'h6bb, 16'h9c70, 16'h9c4f, 16'h9c4f, 16'h94d, 16'h732a, 16'h6aa9, 16'h7b4a, 16'h7b9, 16'h6288, 16'h18a1, 16'h840, 16'h841, 16'h213, 16'h39a5, 16'h39c6, 16'h39a5, 16'h39a5, 16'h39a5, 16'h39a5, 16'h3985, 16'h39a4, 16'h4183, 16'h1881, 16'h840, 16'h840, 16'h840, 16'h840, 16'h840, 16'h1040, 16'h1061, 16'h1061, 16'h1061, 16'h1861, 16'h28e2, 16'h312, 16'h28c1, 16'h49a4, 16'h49e5, 16'h3963, 16'h840, 16'h020, 16'h020, 16'h861, 16'h3165, 16'h5aaa, 16'h6bb, 16'h6bb, 16'h6bb, 16'h6bb, 16'h6bb, 16'h6bb, 16'h6ba, 16'h6aeb, 16'h6bb, 16'h6b2b, 16'h6b2c, 16'h736c, 16'h7bad, 16'h83ae, 16'h83ae, 16'h83ae, 16'h7bad, 16'h7b8d, 16'h7b8d, 16'h7bad, 16'h83ae, 16'h83ae, 16'h83ce, 16'h83ce, 16'h83ce, 16'h83ce, 16'h83ae, 16'h7bad, 16'h7b8d, 16'h7b8d, 16'h734c, 16'h6b2b, 16'h6b2c, 16'h6b2c, 16'h6b2b, 16'h6bb, 16'h6bb, 16'h6bb, 16'h6b2c, 16'h732c, 16'h734c, 16'h7b6d, 16'h9c50, 16'hc574, 16'hc574, 16'hc574, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc553, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb0, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha470, 16'ha470, 16'ha46f, 16'ha46f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h8bac, 16'h41a5, 16'h20e2, 16'h20c2, 16'h20c2, 16'h20c2, 16'h18a1, 16'h820, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'hbd34, 16'hbd13, 16'hbd34, 16'hb514, 16'hb514, 16'hb534, 16'hb533, 16'had13, 16'had13, 16'had13, 16'hacf3, 16'hacf3, 16'hacf3, 16'hacf3, 16'hacf2, 16'ha4d2, 16'h9c70, 16'h8bee, 16'h732b, 16'h3986, 16'h3124, 16'h213, 16'h18c2, 16'h18a2, 16'h18c3, 16'h7b6d, 16'ha4b1, 16'h942f, 16'h8bcd, 16'h8bac, 16'h739, 16'h5a27, 16'h6a88, 16'h6267, 16'h49a5, 16'h1881, 16'h841, 16'h1061, 16'h213, 16'h39c6, 16'h41e6, 16'h427, 16'h4a7, 16'h4a7, 16'h4a7, 16'h49e7, 16'h49e6, 16'h4184, 16'h1061, 16'h020, 16'h020, 16'h020, 16'h020, 16'h820, 16'h820, 16'h1081, 16'h1881, 16'h18a1, 16'h18a1, 16'h3122, 16'h3122, 16'h28e2, 16'h49e4, 16'h51e5, 16'h4184, 16'h1061, 16'h840, 16'h020, 16'h861, 16'h3185, 16'h5aaa, 16'h6bb, 16'h6bb, 16'h6bb, 16'h6bb, 16'h6bb, 16'h6bb, 16'h6bb, 16'h6aeb, 16'h6bb, 16'h6b2b, 16'h732c, 16'h736d, 16'h7bad, 16'h83ae, 16'h83ae, 16'h83ae, 16'h7bad, 16'h7b8d, 16'h7bad, 16'h83ae, 16'h83ce, 16'h83ce, 16'h83ce, 16'h83ae, 16'h83ce, 16'h83ce, 16'h83ae, 16'h7bad, 16'h7b8d, 16'h7b6d, 16'h734c, 16'h6b2b, 16'h6b2b, 16'h6b2b, 16'h6b2b, 16'h6b2c, 16'h6b2c, 16'h734c, 16'h732c, 16'h734c, 16'h734c, 16'h7b6d, 16'h9c50, 16'hc574, 16'hc574, 16'hc574, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc553, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hbd32, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4d2, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h8b8c, 16'h41a5, 16'h20e2, 16'h20c2, 16'h20c2, 16'h20c1, 16'h1881, 16'h820, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'hbcd3, 16'hbcd3, 16'hb534, 16'hb513, 16'hb4f3, 16'hb514, 16'hb533, 16'hb513, 16'had13, 16'had13, 16'hacf3, 16'hacf3, 16'hacf3, 16'hacf3, 16'hacf2, 16'h83ae, 16'h3986, 16'h5248, 16'h6aeb, 16'h20e3, 16'h2925, 16'h20e3, 16'h1061, 16'h861, 16'h1061, 16'h5a89, 16'h9cb1, 16'h942f, 16'h942f, 16'h944f, 16'h7b4b, 16'h49e6, 16'h5a6, 16'h49c5, 16'h20e2, 16'h1881, 16'h18c2, 16'h213, 16'h2924, 16'h39c6, 16'h41e6, 16'h4a7, 16'h4a7, 16'h4a7, 16'h4a7, 16'h4a7, 16'h49e6, 16'h49a4, 16'h20e2, 16'h18a1, 16'h1081, 16'h1081, 16'h1061, 16'h1061, 16'h841, 16'h840, 16'h840, 16'h840, 16'h840, 16'h3122, 16'h3143, 16'h312, 16'h525, 16'h51e5, 16'h4184, 16'h1081, 16'h840, 16'h820, 16'h861, 16'h3165, 16'h5aaa, 16'h6bb, 16'h6b2b, 16'h6b2b, 16'h6b2b, 16'h6b2b, 16'h6b2b, 16'h6bb, 16'h6bb, 16'h6bb, 16'h6b2c, 16'h734c, 16'h7b6d, 16'h7b8d, 16'h7bad, 16'h83ad, 16'h83ad, 16'h7bad, 16'h7b8d, 16'h7bae, 16'h83ce, 16'h83ae, 16'h83ae, 16'h83ae, 16'h83ae, 16'h83ce, 16'h83ce, 16'h7bad, 16'h7bad, 16'h7b8d, 16'h7b6d, 16'h734c, 16'h6b2b, 16'h6b2c, 16'h6b2c, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h6b2c, 16'h734c, 16'h736c, 16'h7b6c, 16'h9c50, 16'hc573, 16'hc574, 16'hc574, 16'hc574, 16'hc573, 16'hc573, 16'hc573, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hbd12, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha46f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h838c, 16'h41a5, 16'h20e2, 16'h20c2, 16'h20c2, 16'h20c1, 16'h1881, 16'h820, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'hb4f3, 16'hb4f3, 16'hb534, 16'hb513, 16'hb4b2, 16'hb4d2, 16'hb534, 16'hb513, 16'had13, 16'had13, 16'had13, 16'had13, 16'hacf3, 16'hacf3, 16'hacf2, 16'h9c91, 16'h83ae, 16'h83ae, 16'h8cf, 16'h39a6, 16'h18c3, 16'h18c2, 16'h10a2, 16'h1061, 16'h1062, 16'h4a8, 16'h9c90, 16'ha4b1, 16'h9c91, 16'h9c90, 16'h8ce, 16'h49e6, 16'h5a6, 16'h49c5, 16'h293, 16'h18a2, 16'h1081, 16'h1881, 16'h213, 16'h39a6, 16'h41e6, 16'h4a7, 16'h4a27, 16'h4a27, 16'h4a27, 16'h4a7, 16'h4a6, 16'h49a4, 16'h20e2, 16'h18a1, 16'h18a2, 16'h18a2, 16'h18c2, 16'h18c2, 16'h18a1, 16'h1061, 16'h860, 16'h820, 16'h820, 16'h3123, 16'h4184, 16'h3963, 16'h5a26, 16'h525, 16'h4184, 16'h1082, 16'h841, 16'h020, 16'h861, 16'h2965, 16'h5aa9, 16'h6bb, 16'h6b2b, 16'h6b2b, 16'h6b2b, 16'h6b2b, 16'h6b2b, 16'h6bb, 16'h6bb, 16'h6bb, 16'h6b2c, 16'h734c, 16'h7b6d, 16'h7bad, 16'h83ae, 16'h83ae, 16'h7bad, 16'h7bad, 16'h7bad, 16'h7bae, 16'h83ae, 16'h83ae, 16'h83ae, 16'h7bae, 16'h83ae, 16'h83ce, 16'h83ce, 16'h7bae, 16'h7b8d, 16'h7b8d, 16'h736d, 16'h732c, 16'h732c, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h736c, 16'h7b6d, 16'h9c70, 16'hc574, 16'hc574, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hbd12, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha470, 16'ha46f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9ce, 16'h838c, 16'h41a5, 16'h20e2, 16'h20c2, 16'h20c2, 16'h20c2, 16'h1881, 16'h820, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'hb554, 16'hb554, 16'hb554, 16'hb534, 16'hb513, 16'hb4f3, 16'hb534, 16'hb534, 16'had13, 16'had13, 16'had13, 16'had13, 16'had13, 16'hacf3, 16'hacf2, 16'hacf2, 16'hacd2, 16'ha4d2, 16'h9450, 16'h6aeb, 16'h39c6, 16'h18c2, 16'h1082, 16'h18a2, 16'h3165, 16'h6b2c, 16'h9cb1, 16'h9cb1, 16'ha4b1, 16'ha4b1, 16'h942e, 16'h41a5, 16'h51e5, 16'h5226, 16'h41a4, 16'h20e2, 16'h1082, 16'h1881, 16'h213, 16'h39a5, 16'h41e6, 16'h4a7, 16'h4a7, 16'h4a27, 16'h4a27, 16'h4a27, 16'h4a6, 16'h49c4, 16'h20e2, 16'h1081, 16'h1061, 16'h841, 16'h861, 16'h1081, 16'h841, 16'h861, 16'h840, 16'h020, 16'h820, 16'h3143, 16'h49a4, 16'h49c5, 16'h5a46, 16'h525, 16'h41a4, 16'h1882, 16'h841, 16'h040, 16'h861, 16'h3185, 16'h5aa9, 16'h6bb, 16'h6b2b, 16'h6b2b, 16'h6b2b, 16'h6b2b, 16'h6b2b, 16'h6b2b, 16'h6bb, 16'h6b2b, 16'h6b2c, 16'h734c, 16'h7b6d, 16'h83ae, 16'h83ae, 16'h83ae, 16'h7bad, 16'h7bad, 16'h7bad, 16'h7bad, 16'h7bad, 16'h7bae, 16'h7bae, 16'h7bae, 16'h7bae, 16'h83ad, 16'h7bad, 16'h7bad, 16'h736d, 16'h6b2d, 16'h62ec, 16'h6bb, 16'h734d, 16'h734c, 16'h734c, 16'h736c, 16'h734c, 16'h734d, 16'h734d, 16'h734c, 16'h734c, 16'h736c, 16'h7b6d, 16'h9c50, 16'hc574, 16'hc574, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb0, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha470, 16'ha44f, 16'ha44f, 16'ha450, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h838c, 16'h4185, 16'h20e2, 16'h20c2, 16'h20c2, 16'h20c2, 16'h1881, 16'h820, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'hb554, 16'hb554, 16'hb554, 16'hb534, 16'hb534, 16'hb534, 16'hb534, 16'hb534, 16'had13, 16'had13, 16'had13, 16'had13, 16'had13, 16'hacf3, 16'hacf3, 16'hacf2, 16'hacf2, 16'hacd2, 16'ha4d2, 16'hacf2, 16'h9470, 16'h4a27, 16'h2924, 16'h427, 16'h7b8d, 16'h9c70, 16'h8ce, 16'h83cd, 16'h8bed, 16'h8ce, 16'h7b8c, 16'h41a5, 16'h51e6, 16'h5a26, 16'h49c4, 16'h2923, 16'h18a2, 16'h18a1, 16'h213, 16'h39a5, 16'h41c6, 16'h49e6, 16'h4a7, 16'h4a7, 16'h4a7, 16'h4a7, 16'h4a6, 16'h49e4, 16'h3983, 16'h2943, 16'h2943, 16'h2123, 16'h2923, 16'h3164, 16'h18a2, 16'h18c3, 16'h10a2, 16'h840, 16'h840, 16'h4184, 16'h526, 16'h5a26, 16'h6246, 16'h525, 16'h41a4, 16'h18a1, 16'h841, 16'h040, 16'h861, 16'h3185, 16'h5aaa, 16'h6bb, 16'h6b2b, 16'h6b2b, 16'h6b2b, 16'h6b2b, 16'h6b2c, 16'h6b2c, 16'h6b2b, 16'h6b2b, 16'h734c, 16'h734c, 16'h7b6d, 16'h83ae, 16'h83ae, 16'h83ce, 16'h7bad, 16'h7bad, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h7bae, 16'h7bae, 16'h7bae, 16'h7bad, 16'h7b8d, 16'h736d, 16'h6b2c, 16'h62ec, 16'h5acb, 16'h5acb, 16'h63b, 16'h736d, 16'h736d, 16'h734c, 16'h734d, 16'h734d, 16'h734c, 16'h736d, 16'h736d, 16'h734c, 16'h736d, 16'h7b8d, 16'h9c50, 16'hc574, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha46f, 16'ha470, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h838c, 16'h4185, 16'h20e2, 16'h20c2, 16'h20c2, 16'h20c2, 16'h1881, 16'h820, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'ha4b2, 16'ha4b2, 16'ha4b2, 16'ha4b2, 16'ha4b2, 16'ha4b2, 16'ha4b2, 16'ha4b2, 16'ha4b2, 16'ha4b2, 16'ha492, 16'ha491, 16'ha491, 16'ha491, 16'ha491, 16'ha491, 16'ha491, 16'ha491, 16'ha4b1, 16'ha4d2, 16'h9470, 16'h5a89, 16'h5268, 16'h7b6c, 16'h942f, 16'h7b8c, 16'h5a88, 16'h5a87, 16'h5a67, 16'h5a88, 16'h5a67, 16'h4a6, 16'h5a26, 16'h5a46, 16'h49c4, 16'h293, 16'h1882, 16'h2944, 16'h213, 16'h39a5, 16'h41c6, 16'h41e6, 16'h4a6, 16'h4a7, 16'h4a7, 16'h4a7, 16'h4a6, 16'h49c4, 16'h20e2, 16'h10a1, 16'h18a1, 16'h18c2, 16'h2123, 16'h4a6, 16'h3985, 16'h2944, 16'h18e3, 16'h861, 16'h840, 16'h4184, 16'h5a26, 16'h5a26, 16'h6266, 16'h5a6, 16'h41a4, 16'h18c2, 16'h861, 16'h840, 16'h881, 16'h3185, 16'h5ac9, 16'h6b2b, 16'h6b2b, 16'h6b2b, 16'h6b2b, 16'h6b2b, 16'h734c, 16'h734c, 16'h6b2c, 16'h734c, 16'h732c, 16'h734c, 16'h7b6d, 16'h7bad, 16'h83ae, 16'h83ad, 16'h7bad, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h7bad, 16'h7b8d, 16'h7b8d, 16'h736d, 16'h6b2c, 16'h62ec, 16'h62ec, 16'h5aeb, 16'h5acb, 16'h5acb, 16'h63b, 16'h736d, 16'h736c, 16'h736d, 16'h734d, 16'h736d, 16'h736d, 16'h736d, 16'h736d, 16'h736d, 16'h736d, 16'h7b6d, 16'h9c4f, 16'hc573, 16'hc574, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc553, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha44f, 16'ha46f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9ce, 16'h836c, 16'h4185, 16'h20e2, 16'h20c2, 16'h20c2, 16'h20c2, 16'h1881, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'hacf3, 16'hacf3, 16'hacf3, 16'ha4d2, 16'ha4d2, 16'ha4b2, 16'ha4b2, 16'ha491, 16'h9c91, 16'h9c71, 16'h9c51, 16'h9450, 16'h9430, 16'h9430, 16'h8cf, 16'h8bef, 16'h8bef, 16'h8bef, 16'h8bce, 16'h83ce, 16'h83ad, 16'h734c, 16'h8bef, 16'h944f, 16'h9c6f, 16'h83cd, 16'h5a88, 16'h5267, 16'h5a67, 16'h6288, 16'h5a47, 16'h5227, 16'h5a47, 16'h5a66, 16'h49c4, 16'h3144, 16'h5228, 16'h734c, 16'h41c6, 16'h3985, 16'h39a5, 16'h41c6, 16'h41e6, 16'h49e6, 16'h4a6, 16'h49e6, 16'h4a6, 16'h49c4, 16'h20c1, 16'h1061, 16'h1061, 16'h1081, 16'h18c2, 16'h41e5, 16'h41c5, 16'h18a2, 16'h020, 16'h020, 16'h840, 16'h4164, 16'h5a26, 16'h5a46, 16'h6a87, 16'h5a26, 16'h49c4, 16'h18c2, 16'h861, 16'h841, 16'h1081, 16'h3185, 16'h5ac9, 16'h6b2b, 16'h6b2b, 16'h6b2b, 16'h6b4b, 16'h6b4c, 16'h734c, 16'h734c, 16'h6b2b, 16'h734c, 16'h734c, 16'h734c, 16'h736d, 16'h7bad, 16'h7bad, 16'h7bad, 16'h7bad, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h736c, 16'h6bc, 16'h62eb, 16'h62eb, 16'h62eb, 16'h5aeb, 16'h62eb, 16'h5acb, 16'h63c, 16'h736d, 16'h7b8d, 16'h736d, 16'h736d, 16'h736d, 16'h736d, 16'h736d, 16'h736d, 16'h736d, 16'h736c, 16'h7b6d, 16'h9c4f, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc553, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd52, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9ce, 16'h836c, 16'h4185, 16'h20e2, 16'h20e2, 16'h20c2, 16'h20c1, 16'h1881, 16'h820, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'hb554, 16'hb554, 16'hb534, 16'hb534, 16'hb534, 16'hb534, 16'hb533, 16'had13, 16'had13, 16'had13, 16'hacf3, 16'hacf3, 16'hacf3, 16'hacf2, 16'ha4d2, 16'ha4d2, 16'ha4d2, 16'ha4b2, 16'ha4b2, 16'ha491, 16'h9c91, 16'h9c91, 16'h9c71, 16'h9c90, 16'h9c90, 16'h8bee, 16'h62a8, 16'h5a67, 16'h5a67, 16'h6288, 16'h5a67, 16'h527, 16'h5a48, 16'h6287, 16'h49c5, 16'h49c5, 16'h6aea, 16'h734b, 16'h4a6, 16'h3164, 16'h3164, 16'h3984, 16'h3985, 16'h39a5, 16'h39a5, 16'h3985, 16'h49c5, 16'h49e4, 16'h3143, 16'h213, 16'h213, 16'h213, 16'h20e2, 16'h39a5, 16'h41e5, 16'h18c2, 16'h841, 16'h840, 16'h841, 16'h4184, 16'h6267, 16'h6aa8, 16'h7ae9, 16'h5a46, 16'h49c4, 16'h20c2, 16'h1081, 16'h861, 16'h1081, 16'h3165, 16'h5aa9, 16'h6b2b, 16'h6b4b, 16'h6b2b, 16'h6b4c, 16'h6b4c, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h736d, 16'h7b8d, 16'h7b8d, 16'h7bad, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h7b6d, 16'h7b8d, 16'h7b8d, 16'h736d, 16'h734c, 16'h63b, 16'h63b, 16'h62eb, 16'h62eb, 16'h62ec, 16'h62ec, 16'h5acc, 16'h6bc, 16'h7b8d, 16'h7b8d, 16'h7b6d, 16'h7b6d, 16'h736d, 16'h736d, 16'h736d, 16'h7b6d, 16'h736d, 16'h736d, 16'h7b6d, 16'h9c50, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc553, 16'hc553, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'hac90, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha470, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha450, 16'ha450, 16'ha450, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9ce, 16'h836c, 16'h3984, 16'h20e2, 16'h20c1, 16'h20c2, 16'h20c2, 16'h1081, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'hb554, 16'hb554, 16'hb554, 16'hb534, 16'hb534, 16'hb534, 16'hb534, 16'hb513, 16'hb513, 16'had13, 16'had13, 16'had13, 16'hacf3, 16'hacf2, 16'hacf2, 16'ha4d2, 16'ha4d2, 16'ha4d2, 16'ha4d2, 16'ha4b2, 16'ha4b1, 16'ha4b1, 16'ha491, 16'ha490, 16'h9c90, 16'h8bee, 16'h5a88, 16'h5a87, 16'h4a26, 16'h5a67, 16'h62a8, 16'h5247, 16'h6aa9, 16'h6287, 16'h49e4, 16'h49e5, 16'h525, 16'h525, 16'h49e5, 16'h525, 16'h525, 16'h51e5, 16'h51e5, 16'h51e5, 16'h49e5, 16'h49c4, 16'h51e4, 16'h51e4, 16'h49c4, 16'h49a4, 16'h49a4, 16'h41a4, 16'h41a4, 16'h49c5, 16'h49e5, 16'h41a4, 16'h3984, 16'h3143, 16'h3123, 16'h49c4, 16'h5a46, 16'h6267, 16'h6a87, 16'h5a25, 16'h49c4, 16'h2923, 16'h213, 16'h18c2, 16'h1082, 16'h214, 16'h5aa9, 16'h6b4b, 16'h6b4b, 16'h6b2b, 16'h6b2c, 16'h6b4c, 16'h6b2c, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h736c, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h7b6d, 16'h736d, 16'h736d, 16'h736d, 16'h7b8d, 16'h7b8d, 16'h736d, 16'h734d, 16'h63c, 16'h63c, 16'h62ec, 16'h62eb, 16'h62ec, 16'h62ec, 16'h62ec, 16'h6b2c, 16'h7b8d, 16'h7b8d, 16'h7b6d, 16'h7b6d, 16'h736d, 16'h736d, 16'h736d, 16'h736d, 16'h736d, 16'h7b6d, 16'h7b6d, 16'h9c50, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc553, 16'hc553, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacd1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'hac90, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha46f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9ce, 16'h836c, 16'h3984, 16'h20e2, 16'h20c2, 16'h20c2, 16'h20c2, 16'h1081, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'hb554, 16'hb554, 16'hb554, 16'hb554, 16'hb534, 16'hb534, 16'hb534, 16'hb534, 16'hb534, 16'hb514, 16'hb513, 16'hb534, 16'hacf3, 16'h9c91, 16'ha4b2, 16'ha4b2, 16'ha4b2, 16'ha4b2, 16'ha4d2, 16'ha4b2, 16'ha4b1, 16'ha4b1, 16'ha491, 16'h9c90, 16'ha490, 16'h8bed, 16'h5a87, 16'h5226, 16'h39a4, 16'h41c5, 16'h4a6, 16'h49e5, 16'h6ae9, 16'h5226, 16'h49e5, 16'h4a6, 16'h20e3, 16'h20e2, 16'h3143, 16'h62a9, 16'h6aea, 16'h6ac9, 16'h6aea, 16'h6ac9, 16'h51e5, 16'h49a4, 16'h525, 16'h51e5, 16'h49e4, 16'h49a4, 16'h49a4, 16'h49c4, 16'h49c4, 16'h525, 16'h525, 16'h5226, 16'h525, 16'h49c4, 16'h49c4, 16'h525, 16'h5a26, 16'h5a26, 16'h5a25, 16'h525, 16'h5226, 16'h4a26, 16'h3184, 16'h2944, 16'h20e2, 16'h2924, 16'h5ac9, 16'h6b4b, 16'h6b2b, 16'h6b2b, 16'h6b2b, 16'h6b2b, 16'h6b2c, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h736c, 16'h7b8d, 16'h7b6d, 16'h7b6d, 16'h736d, 16'h736d, 16'h736d, 16'h7b6d, 16'h7b8d, 16'h7b6d, 16'h736d, 16'h736d, 16'h63c, 16'h63c, 16'h63c, 16'h63c, 16'h63c, 16'h62ec, 16'h62ec, 16'h6b2c, 16'h738d, 16'h7b8d, 16'h736d, 16'h736d, 16'h736d, 16'h736d, 16'h734d, 16'h736d, 16'h736d, 16'h7b6d, 16'h7b6d, 16'h9c50, 16'hc573, 16'hc574, 16'hc574, 16'hc573, 16'hc573, 16'hc573, 16'hc553, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'ha490, 16'ha490, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha470, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h94e, 16'h836b, 16'h3984, 16'h20e2, 16'h20c2, 16'h20c2, 16'h20c2, 16'h1081, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'hbd54, 16'hb554, 16'hb534, 16'hb554, 16'hb534, 16'hb534, 16'hb534, 16'hb534, 16'hb534, 16'hb514, 16'hacf3, 16'hacf3, 16'hacf3, 16'h9451, 16'ha4b2, 16'ha4b2, 16'ha492, 16'ha4b1, 16'ha4d2, 16'ha4b2, 16'ha4b2, 16'ha4b1, 16'h8bef, 16'h8bcd, 16'ha490, 16'h8bed, 16'h5a67, 16'h39a4, 16'h18e2, 16'h18e2, 16'h18e2, 16'h2923, 16'h4a5, 16'h3984, 16'h293, 16'h293, 16'h1861, 16'h1881, 16'h1881, 16'h3144, 16'h3144, 16'h3964, 16'h41a5, 16'h3964, 16'h28e2, 16'h28e2, 16'h49a4, 16'h4183, 16'h292, 16'h20c1, 16'h20e2, 16'h28e2, 16'h20e2, 16'h3143, 16'h3963, 16'h3984, 16'h3143, 16'h20c2, 16'h20a1, 16'h4184, 16'h6267, 16'h5a26, 16'h41a4, 16'h3143, 16'h2923, 16'h2964, 16'h2944, 16'h39a5, 16'h39a5, 16'h4a27, 16'h6ba, 16'h6b4c, 16'h6b2c, 16'h6b2b, 16'h6b2b, 16'h6b2c, 16'h6b2c, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h7b6d, 16'h7b6d, 16'h7b8d, 16'h736d, 16'h736c, 16'h7b6c, 16'h7b6d, 16'h7b6d, 16'h7b6d, 16'h736d, 16'h736c, 16'h6b2c, 16'h63c, 16'h63c, 16'h62ec, 16'h62ec, 16'h62ec, 16'h62ec, 16'h6b2c, 16'h7b8d, 16'h736d, 16'h736d, 16'h736d, 16'h736d, 16'h736d, 16'h736d, 16'h736d, 16'h736c, 16'h736c, 16'h7b6d, 16'ha470, 16'hc573, 16'hc574, 16'hc574, 16'hc573, 16'hc573, 16'hc573, 16'hc553, 16'hc553, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hbd12, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9ce, 16'h94e, 16'h836c, 16'h3984, 16'h20e2, 16'h20c2, 16'h20c2, 16'h20c2, 16'h1081, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'hb554, 16'hb533, 16'hacf3, 16'hb534, 16'hb513, 16'had13, 16'hb534, 16'hb534, 16'hb534, 16'hacf3, 16'hacd3, 16'hacf3, 16'hacd3, 16'h9430, 16'ha492, 16'ha4b2, 16'ha4b2, 16'ha491, 16'ha4d2, 16'ha4b2, 16'ha4b1, 16'ha4b1, 16'h8bee, 16'h838c, 16'ha490, 16'h83ad, 16'h5a47, 16'h39a5, 16'h213, 16'h213, 16'h193, 16'h213, 16'h39a4, 16'h732a, 16'h7b4a, 16'h5a88, 16'h3965, 16'h20e3, 16'h2924, 16'h5268, 16'h62ea, 16'h6ba, 16'h6aea, 16'h62a9, 16'h5248, 16'h41a5, 16'h3984, 16'h2923, 16'h20e2, 16'h20e2, 16'h20e2, 16'h20e2, 16'h212, 16'h3984, 16'h3964, 16'h3964, 16'h3123, 16'h20c2, 16'h20c2, 16'h3143, 16'h5226, 16'h41c5, 16'h2923, 16'h20e2, 16'h1081, 16'h1061, 16'h20e3, 16'h41c6, 16'h427, 16'h5288, 16'h6bb, 16'h6b2c, 16'h6b2c, 16'h6b2b, 16'h6b2b, 16'h6b2c, 16'h732c, 16'h734c, 16'h734c, 16'h734c, 16'h732c, 16'h6b2c, 16'h6b2c, 16'h736c, 16'h7b6c, 16'h7b8d, 16'h736d, 16'h736d, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h7b6d, 16'h736d, 16'h6b2c, 16'h6bc, 16'h63c, 16'h62ec, 16'h63c, 16'h63c, 16'h63c, 16'h6bc, 16'h736d, 16'h736d, 16'h736d, 16'h736d, 16'h736d, 16'h736d, 16'h736c, 16'h736c, 16'h736c, 16'h736c, 16'h7b6d, 16'ha470, 16'hc573, 16'hc574, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc553, 16'hc553, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd52, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hbd12, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9ce, 16'h9ce, 16'h836c, 16'h3984, 16'h20e2, 16'h20c2, 16'h20c2, 16'h18c2, 16'h1081, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'hacf2, 16'hacf3, 16'hacf3, 16'hacf3, 16'hb513, 16'hb513, 16'hb534, 16'hb534, 16'hb534, 16'hacf3, 16'hacd3, 16'hacd3, 16'hacd3, 16'h9450, 16'h9c72, 16'ha492, 16'ha4b2, 16'ha4b2, 16'ha4d2, 16'ha4b2, 16'ha4b2, 16'ha4b1, 16'h9c70, 16'h83ad, 16'h8bee, 16'h83cd, 16'h5247, 16'h39c5, 16'h213, 16'h2123, 16'h2123, 16'h2123, 16'h39a4, 16'h62c9, 16'h83ac, 16'h83ad, 16'h83ad, 16'h736c, 16'h5a69, 16'h41a6, 16'h3985, 16'h4a7, 16'h62ca, 16'h62ea, 16'h5aa9, 16'h41e6, 16'h3164, 16'h213, 16'h213, 16'h213, 16'h2923, 16'h2943, 16'h2943, 16'h5a68, 16'h5247, 16'h4a27, 16'h3985, 16'h18a2, 16'h1061, 16'h213, 16'h427, 16'h3184, 16'h18e2, 16'h2923, 16'h293, 16'h18c2, 16'h2924, 16'h4a7, 16'h5268, 16'h5aa9, 16'h6bb, 16'h6b2c, 16'h6b4c, 16'h6b2c, 16'h6b2c, 16'h6b2c, 16'h6b4c, 16'h734c, 16'h734c, 16'h6b4c, 16'h6b2c, 16'h6b2c, 16'h6b4c, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h7b6d, 16'h7b6d, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h736d, 16'h6b2c, 16'h6b2c, 16'h63c, 16'h63c, 16'h63c, 16'h62ec, 16'h62ec, 16'h6bc, 16'h736d, 16'h736d, 16'h736d, 16'h736c, 16'h736d, 16'h736d, 16'h736d, 16'h736c, 16'h736c, 16'h736c, 16'h7b6c, 16'h9c4f, 16'hc573, 16'hc574, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc553, 16'hc553, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hbd12, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9ce, 16'h94e, 16'h836c, 16'h3964, 16'h20c2, 16'h20c2, 16'h20c2, 16'h20c1, 16'h1081, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'hacf2, 16'hacf3, 16'hacf3, 16'hacf3, 16'hb534, 16'hb514, 16'hb534, 16'hb534, 16'hb534, 16'hb534, 16'hb514, 16'hacf3, 16'hacf3, 16'h9c92, 16'ha492, 16'ha492, 16'ha4b2, 16'ha4d2, 16'ha4d2, 16'ha4b2, 16'ha4b2, 16'ha4b1, 16'h9c91, 16'h942f, 16'h838c, 16'h7b6c, 16'h5a67, 16'h39a5, 16'h193, 16'h2123, 16'h2123, 16'h2123, 16'h3184, 16'h2923, 16'h62a9, 16'h732b, 16'h734c, 16'h734c, 16'h734c, 16'h6bb, 16'h5269, 16'h3186, 16'h214, 16'h213, 16'h20e4, 16'h18c2, 16'h18c2, 16'h18c2, 16'h212, 16'h2923, 16'h2923, 16'h2923, 16'h3143, 16'h5a88, 16'h5267, 16'h4a47, 16'h31a5, 16'h10a2, 16'h1061, 16'h18e2, 16'h41e6, 16'h2944, 16'h10a2, 16'h10a2, 16'h18c2, 16'h20e2, 16'h3164, 16'h5289, 16'h62ca, 16'h62ea, 16'h6b2b, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h6b4c, 16'h734c, 16'h734c, 16'h6b2c, 16'h6b4c, 16'h734c, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h738d, 16'h6b2c, 16'h63c, 16'h63c, 16'h63c, 16'h63c, 16'h62ec, 16'h62ec, 16'h6b2c, 16'h7b6d, 16'h736d, 16'h736d, 16'h736c, 16'h736d, 16'h736d, 16'h736d, 16'h736c, 16'h736c, 16'h736c, 16'h7b6c, 16'h9c4f, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc553, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd52, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd0, 16'hacb0, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha44f, 16'ha46f, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h94e, 16'h7b6b, 16'h3964, 16'h20e2, 16'h20c2, 16'h20c2, 16'h20c1, 16'h1881, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'hb534, 16'hb513, 16'hacf3, 16'hb534, 16'hb534, 16'hb534, 16'hb534, 16'hb534, 16'hb534, 16'hb513, 16'ha4d2, 16'hacd2, 16'hacf3, 16'hacf3, 16'hacf3, 16'hacf2, 16'hacd2, 16'ha4d2, 16'ha4d2, 16'ha4d2, 16'ha4b2, 16'ha4b1, 16'h9c91, 16'h942f, 16'h734b, 16'h734b, 16'h5a67, 16'h39a5, 16'h212, 16'h212, 16'h2123, 16'h213, 16'h3184, 16'h293, 16'h5a89, 16'h734c, 16'h7b6d, 16'h7b6d, 16'h7b6d, 16'h7b6d, 16'h734c, 16'h734c, 16'h62ea, 16'h41c7, 16'h20c3, 16'h1082, 16'h10a2, 16'h1081, 16'h1061, 16'h1081, 16'h1081, 16'h1081, 16'h293, 16'h62a8, 16'h5a67, 16'h4a48, 16'h39a6, 16'h1882, 16'h861, 16'h18a2, 16'h39c6, 16'h2944, 16'h10a2, 16'h1082, 16'h18a2, 16'h18c2, 16'h3164, 16'h5aa9, 16'h62eb, 16'h6b2b, 16'h734c, 16'h734c, 16'h736c, 16'h736c, 16'h736c, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h7b6d, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h736d, 16'h736d, 16'h6b2c, 16'h63c, 16'h63c, 16'h63b, 16'h62ec, 16'h62ec, 16'h62ec, 16'h6bc, 16'h7b8d, 16'h736d, 16'h736d, 16'h736d, 16'h736d, 16'h736d, 16'h736d, 16'h736c, 16'h736c, 16'h7b6c, 16'h7b6d, 16'h9c4f, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc553, 16'hc553, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9ce, 16'h834b, 16'h3964, 16'h20e2, 16'h20c2, 16'h20c2, 16'h20c2, 16'h1081, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'hb554, 16'hb534, 16'hb534, 16'hb534, 16'hb534, 16'hb534, 16'hb534, 16'hb554, 16'hacd2, 16'h9c71, 16'ha492, 16'ha492, 16'h9c91, 16'hacf2, 16'hacf3, 16'hacf2, 16'hacf2, 16'ha4d2, 16'ha4d2, 16'ha4b2, 16'ha4b2, 16'ha4b1, 16'h9cb1, 16'h9c70, 16'h734c, 16'h5a88, 16'h5226, 16'h5247, 16'h4a6, 16'h4a6, 16'h4a6, 16'h4a6, 16'h39a5, 16'h20c2, 16'h5a89, 16'h7b6c, 16'h83ad, 16'h83ad, 16'h83ad, 16'h83ad, 16'h83ad, 16'h83ad, 16'h83ad, 16'h6bb, 16'h5248, 16'h41e6, 16'h41c6, 16'h3165, 16'h18c3, 16'h1081, 16'h861, 16'h861, 16'h2923, 16'h6ac9, 16'h5267, 16'h4a47, 16'h3164, 16'h1081, 16'h840, 16'h841, 16'h3185, 16'h2124, 16'h861, 16'h1081, 16'h18a2, 16'h18c2, 16'h3185, 16'h62ea, 16'h6b2b, 16'h6b4c, 16'h734c, 16'h734c, 16'h734c, 16'h736c, 16'h736c, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h736d, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h7b6d, 16'h7b6d, 16'h736d, 16'h6b2c, 16'h63c, 16'h63c, 16'h63c, 16'h62ec, 16'h62ec, 16'h62ec, 16'h6bc, 16'h736d, 16'h7b6d, 16'h736d, 16'h736d, 16'h736d, 16'h736d, 16'h736d, 16'h734c, 16'h734c, 16'h7b6d, 16'h7b6d, 16'h9c4f, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc553, 16'hc553, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha470, 16'ha46f, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9ce, 16'h7b4b, 16'h3964, 16'h20e2, 16'h20c2, 16'h20c2, 16'h20c2, 16'h1081, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'hb554, 16'hb554, 16'hb554, 16'hb554, 16'hb554, 16'hb534, 16'hb534, 16'ha492, 16'h9450, 16'ha4b2, 16'ha4b2, 16'hacd2, 16'ha4d2, 16'ha4b1, 16'ha4b2, 16'hacf2, 16'hacf2, 16'hacd2, 16'ha4d2, 16'ha4d2, 16'ha4d2, 16'ha4b2, 16'h9cb1, 16'h9cb1, 16'h9c91, 16'h7b8d, 16'h5a68, 16'h4a7, 16'h41a5, 16'h49e6, 16'h41e6, 16'h5267, 16'h41c6, 16'h3144, 16'h5227, 16'h5248, 16'h4a7, 16'h5227, 16'h5247, 16'h5248, 16'h5268, 16'h5a88, 16'h62a9, 16'h62a9, 16'h62a9, 16'h62a9, 16'h62a9, 16'h5aa9, 16'h5268, 16'h41c5, 16'h3144, 16'h3144, 16'h41e5, 16'h6ae9, 16'h5247, 16'h39c6, 16'h20e3, 16'h861, 16'h841, 16'h861, 16'h39c6, 16'h2944, 16'h861, 16'h10a2, 16'h213, 16'h39a5, 16'h5268, 16'h6bb, 16'h6b2c, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h736c, 16'h736d, 16'h736c, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h7b6d, 16'h7b8d, 16'h7b8d, 16'h736d, 16'h736d, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h736d, 16'h6b2c, 16'h63c, 16'h63c, 16'h63c, 16'h62ec, 16'h62ec, 16'h62ec, 16'h6b2c, 16'h738d, 16'h736d, 16'h736c, 16'h736d, 16'h736d, 16'h736d, 16'h736c, 16'h736c, 16'h736c, 16'h7b6d, 16'h7b6c, 16'h9c4f, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc553, 16'hc553, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h94e, 16'h836b, 16'h3964, 16'h20c2, 16'h20c2, 16'h20c2, 16'h18c2, 16'h1081, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'hb534, 16'hb554, 16'hb554, 16'hb554, 16'hb554, 16'hb534, 16'h9c71, 16'h9c51, 16'hacf3, 16'hb513, 16'ha4b2, 16'ha4d2, 16'hb513, 16'hacf3, 16'ha4b2, 16'h9c91, 16'ha4d2, 16'hacd2, 16'ha4d2, 16'ha4d2, 16'ha4d2, 16'ha4d2, 16'ha4b2, 16'h9cb1, 16'h9c91, 16'h9c70, 16'h83ae, 16'h5a69, 16'h41a5, 16'h62a9, 16'h6aeb, 16'h732b, 16'h5a89, 16'h5268, 16'h62ca, 16'h6aea, 16'h6aca, 16'h62a9, 16'h6289, 16'h62a9, 16'h62a9, 16'h62c9, 16'h62c9, 16'h62a9, 16'h62a9, 16'h62a9, 16'h5aa9, 16'h5a89, 16'h5a88, 16'h5247, 16'h49e6, 16'h4a27, 16'h5247, 16'h41c5, 16'h213, 16'h1081, 16'h1081, 16'h18e3, 16'h2924, 16'h3185, 16'h5268, 16'h3185, 16'h2944, 16'h4a27, 16'h5aa9, 16'h6b2b, 16'h6b4c, 16'h6b2b, 16'h6b2c, 16'h734c, 16'h734c, 16'h6b2b, 16'h6b2b, 16'h734c, 16'h736d, 16'h736c, 16'h736c, 16'h734c, 16'h734c, 16'h736c, 16'h734c, 16'h734c, 16'h734c, 16'h7b6d, 16'h7b6d, 16'h7b6d, 16'h7b6d, 16'h7b6d, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h736d, 16'h6b2c, 16'h63c, 16'h63c, 16'h63b, 16'h62ec, 16'h62ec, 16'h62ec, 16'h63c, 16'h736c, 16'h736c, 16'h736c, 16'h736d, 16'h736d, 16'h734c, 16'h734c, 16'h736c, 16'h736d, 16'h736d, 16'h7b6d, 16'h9c4f, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc553, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hbd12, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h94e, 16'h834b, 16'h3964, 16'h20c2, 16'h20c2, 16'h20c2, 16'h18c2, 16'h1081, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'hb534, 16'hb554, 16'hb554, 16'hb554, 16'hb554, 16'hb554, 16'hacf3, 16'hb534, 16'hacf3, 16'h9c71, 16'ha4b2, 16'hacd2, 16'hacd2, 16'hacf3, 16'had13, 16'ha4b2, 16'h9c71, 16'hacd2, 16'hacf2, 16'ha4d2, 16'ha4d2, 16'ha4d2, 16'ha4d2, 16'h9cb1, 16'h9c91, 16'h9470, 16'h9450, 16'h8bef, 16'h62ca, 16'h732c, 16'h8bef, 16'h83ce, 16'h83ad, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h732b, 16'h6aca, 16'h7b4d, 16'h7b8d, 16'h7b8d, 16'h7b6d, 16'h7b6d, 16'h7b6d, 16'h7b4c, 16'h734c, 16'h732c, 16'h732c, 16'h5268, 16'h3144, 16'h41e6, 16'h4a28, 16'h2944, 16'h18c2, 16'h214, 16'h2924, 16'h39a5, 16'h427, 16'h4a48, 16'h5289, 16'h5aaa, 16'h6b2b, 16'h734c, 16'h734c, 16'h736c, 16'h734c, 16'h6bc, 16'h6b2c, 16'h734c, 16'h6b4c, 16'h6b2b, 16'h6b2b, 16'h734c, 16'h736d, 16'h736c, 16'h736c, 16'h734c, 16'h736c, 16'h736c, 16'h6b4c, 16'h734c, 16'h734c, 16'h736d, 16'h7b6d, 16'h7b6d, 16'h7b6d, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h738d, 16'h736d, 16'h736d, 16'h6b2c, 16'h63c, 16'h63c, 16'h62ec, 16'h5aec, 16'h62ec, 16'h62ec, 16'h63c, 16'h736c, 16'h736d, 16'h736d, 16'h736d, 16'h736c, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h736c, 16'h7b6d, 16'h9c4f, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc553, 16'hc553, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd52, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h94e, 16'h7b4b, 16'h3964, 16'h20e2, 16'h20c2, 16'h20c2, 16'h20c2, 16'h1081, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'hb554, 16'hb534, 16'hb554, 16'hb554, 16'hb554, 16'hb534, 16'hb554, 16'ha4d2, 16'h9451, 16'ha492, 16'ha4b2, 16'hacd3, 16'hacf3, 16'ha4b2, 16'hacf2, 16'h9c91, 16'h9c71, 16'hacf2, 16'hacf2, 16'hacf2, 16'ha4f2, 16'ha4f2, 16'ha4d2, 16'ha4b1, 16'h9c91, 16'h9c70, 16'h9450, 16'h9430, 16'h8cf, 16'h8cf, 16'h8cf, 16'h8bef, 16'h8bcf, 16'h8bce, 16'h83ce, 16'h83ce, 16'h83ce, 16'h83ae, 16'h838e, 16'h838e, 16'h7b8d, 16'h7b8d, 16'h7b6d, 16'h7b6d, 16'h7b6d, 16'h7b6d, 16'h7b4c, 16'h734c, 16'h734c, 16'h5268, 16'h3144, 16'h41c6, 16'h4a28, 16'h3165, 16'h213, 16'h4a48, 16'h4a48, 16'h4a27, 16'h4a28, 16'h428, 16'h4a49, 16'h6bb, 16'h736d, 16'h736d, 16'h734c, 16'h736c, 16'h734c, 16'h6bb, 16'h6b2c, 16'h734c, 16'h734c, 16'h6b2b, 16'h6b2b, 16'h736c, 16'h736d, 16'h736c, 16'h736c, 16'h734c, 16'h736c, 16'h736d, 16'h734c, 16'h734c, 16'h734c, 16'h736c, 16'h7b8d, 16'h7b8d, 16'h736d, 16'h7b6d, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h738d, 16'h736d, 16'h734c, 16'h6b2c, 16'h63c, 16'h63c, 16'h62eb, 16'h62eb, 16'h5aec, 16'h5aeb, 16'h63c, 16'h736c, 16'h736c, 16'h736d, 16'h736c, 16'h736c, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h736c, 16'h7b6d, 16'h9c2f, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc553, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha46f, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h94e, 16'h7b4b, 16'h3964, 16'h20c2, 16'h20c2, 16'h20c2, 16'h20c2, 16'h1081, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'hb555, 16'hb554, 16'hb554, 16'hb534, 16'hb534, 16'hb554, 16'h9c91, 16'h9451, 16'ha4d3, 16'hacf3, 16'ha4d2, 16'hacd3, 16'hb534, 16'hb513, 16'ha4b2, 16'h9450, 16'hacf2, 16'hacf3, 16'hacf3, 16'hacf3, 16'had13, 16'hacf2, 16'ha4d2, 16'ha4b2, 16'h9c91, 16'h9450, 16'h9430, 16'h8c2f, 16'h7bae, 16'h736d, 16'h736d, 16'h736d, 16'h736c, 16'h734c, 16'h736c, 16'h7b6c, 16'h7b6c, 16'h7b6d, 16'h7b6d, 16'h7b4d, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h732c, 16'h732c, 16'h732b, 16'h5268, 16'h3124, 16'h41c6, 16'h4a28, 16'h2944, 16'h213, 16'h5268, 16'h5268, 16'h5268, 16'h4a48, 16'h428, 16'h4a49, 16'h6bb, 16'h736d, 16'h736d, 16'h734c, 16'h736c, 16'h734c, 16'h6bb, 16'h6b2c, 16'h734c, 16'h734c, 16'h6b2c, 16'h6b2b, 16'h736c, 16'h7b6d, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h736d, 16'h734c, 16'h734c, 16'h6b2b, 16'h736d, 16'h7b6d, 16'h736d, 16'h736d, 16'h736d, 16'h7b6d, 16'h7b8d, 16'h7b8d, 16'h738d, 16'h736d, 16'h736d, 16'h6b2c, 16'h63c, 16'h63b, 16'h62eb, 16'h62eb, 16'h5aeb, 16'h5acc, 16'h63c, 16'h736d, 16'h736d, 16'h736c, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h736c, 16'h7b6d, 16'h9c2f, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc553, 16'hc553, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha470, 16'ha46f, 16'ha46f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9ce, 16'h7b4b, 16'h3964, 16'h20e2, 16'h20c2, 16'h20c2, 16'h20c2, 16'h1081, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'hb534, 16'hb534, 16'hb535, 16'hb535, 16'hb534, 16'hb534, 16'ha4d2, 16'had13, 16'ha492, 16'h9c51, 16'hacf3, 16'hb534, 16'hb514, 16'hb534, 16'hb534, 16'hacf2, 16'h9c91, 16'hacf3, 16'had13, 16'hb534, 16'hb554, 16'hb513, 16'ha4d2, 16'h94f, 16'h9c91, 16'h83ce, 16'h7b6d, 16'h736c, 16'h3985, 16'h18c2, 16'h18c2, 16'h18c2, 16'h18c2, 16'h18c2, 16'h18c3, 16'h20e3, 16'h20e3, 16'h20e3, 16'h213, 16'h213, 16'h213, 16'h214, 16'h2124, 16'h2924, 16'h2924, 16'h2924, 16'h2944, 16'h2944, 16'h2944, 16'h213, 16'h1081, 16'h20e3, 16'h213, 16'h1082, 16'h18c3, 16'h5269, 16'h5a89, 16'h5aaa, 16'h5289, 16'h4a49, 16'h526a, 16'h6b2c, 16'h7b8d, 16'h736d, 16'h734c, 16'h736d, 16'h734c, 16'h6b2c, 16'h6b4c, 16'h736c, 16'h734c, 16'h6b2c, 16'h6b2b, 16'h734c, 16'h736d, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h736c, 16'h734c, 16'h734c, 16'h6b2c, 16'h734c, 16'h736c, 16'h736c, 16'h736c, 16'h736d, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h7b6d, 16'h736d, 16'h736c, 16'h6bc, 16'h63c, 16'h63b, 16'h62ec, 16'h5aeb, 16'h5acb, 16'h5acb, 16'h63c, 16'h736d, 16'h736c, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h734d, 16'h734d, 16'h942f, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc553, 16'hc553, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9cf, 16'h9ce, 16'h94e, 16'h7b4b, 16'h3164, 16'h20e2, 16'h20c2, 16'h20c2, 16'h20c2, 16'h1081, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'had14, 16'hb534, 16'hb514, 16'hb534, 16'hb534, 16'hb554, 16'hb534, 16'h9c71, 16'h9451, 16'hacd3, 16'ha4b2, 16'hacf3, 16'hb534, 16'hb534, 16'hb534, 16'hacf3, 16'h9c91, 16'had13, 16'hb534, 16'hb554, 16'hb553, 16'hb553, 16'hb513, 16'h9c50, 16'h9c70, 16'h83ad, 16'h734b, 16'h6b2b, 16'h20e3, 16'h861, 16'h840, 16'h840, 16'h840, 16'h840, 16'h841, 16'h841, 16'h840, 16'h840, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h840, 16'h840, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h840, 16'h1082, 16'h4a48, 16'h62ca, 16'h62cb, 16'h62cb, 16'h528a, 16'h528a, 16'h6b2c, 16'h736d, 16'h736d, 16'h734c, 16'h736d, 16'h734c, 16'h6b2c, 16'h734c, 16'h736c, 16'h734c, 16'h6b4c, 16'h6b2b, 16'h6b4c, 16'h736c, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h736c, 16'h734c, 16'h734c, 16'h6b2c, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h736d, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h736d, 16'h736c, 16'h6bb, 16'h63b, 16'h63b, 16'h62ec, 16'h5aeb, 16'h5acb, 16'h5aeb, 16'h63c, 16'h734d, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h732c, 16'h732c, 16'h734c, 16'h734c, 16'h942f, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hbd12, 16'hbd12, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9ce, 16'h94e, 16'h7b4b, 16'h3144, 16'h20e2, 16'h20c2, 16'h20c2, 16'h20c2, 16'h1081, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'hacf3, 16'hacf4, 16'h9c71, 16'ha492, 16'hb514, 16'hb534, 16'h9c72, 16'h9c71, 16'hacf3, 16'hb554, 16'hacd3, 16'hb514, 16'hb554, 16'hbd55, 16'hb514, 16'ha4d2, 16'had13, 16'hb554, 16'hb554, 16'hbd75, 16'hb553, 16'hb553, 16'hb553, 16'hacf2, 16'h9c90, 16'h8bee, 16'h8bed, 16'h7b6c, 16'h213, 16'h861, 16'h840, 16'h840, 16'h840, 16'h840, 16'h840, 16'h840, 16'h840, 16'h040, 16'h040, 16'h840, 16'h840, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h020, 16'h020, 16'h020, 16'h040, 16'h840, 16'h840, 16'h840, 16'h1081, 16'h4a48, 16'h62ca, 16'h62eb, 16'h62cb, 16'h528a, 16'h528a, 16'h6b2c, 16'h736d, 16'h736d, 16'h736c, 16'h736c, 16'h734c, 16'h6b2c, 16'h6b4c, 16'h736c, 16'h734c, 16'h6b4c, 16'h6b2c, 16'h6b4c, 16'h736c, 16'h734c, 16'h734c, 16'h734c, 16'h736c, 16'h734c, 16'h734c, 16'h734c, 16'h732c, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h734d, 16'h7b8d, 16'h738d, 16'h736d, 16'h7b6d, 16'h736d, 16'h734d, 16'h6bb, 16'h63b, 16'h62eb, 16'h5aec, 16'h62ec, 16'h62eb, 16'h5aeb, 16'h6bc, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h942f, 16'hc553, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd52, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hbd12, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb0, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h94e, 16'h7b4b, 16'h3944, 16'h20e2, 16'h20e2, 16'h20c2, 16'h20c2, 16'h1081, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'ha4d3, 16'hacf3, 16'ha4b3, 16'ha4d3, 16'had14, 16'hb554, 16'hacf3, 16'hbd55, 16'hbd55, 16'hc595, 16'hbd55, 16'hb534, 16'hb534, 16'hb554, 16'hbd75, 16'hbd75, 16'had13, 16'hb554, 16'hb554, 16'hbd95, 16'had12, 16'h8cf, 16'h8cf, 16'h8bee, 16'h83ad, 16'h83ad, 16'ha4d1, 16'h83ad, 16'h2923, 16'h861, 16'h840, 16'h840, 16'h840, 16'h840, 16'h840, 16'h840, 16'h840, 16'h840, 16'h840, 16'h840, 16'h840, 16'h840, 16'h840, 16'h040, 16'h040, 16'h040, 16'h040, 16'h840, 16'h840, 16'h040, 16'h040, 16'h040, 16'h040, 16'h841, 16'h1081, 16'h4a48, 16'h62cb, 16'h62eb, 16'h62eb, 16'h528a, 16'h528a, 16'h6bc, 16'h736d, 16'h7b6d, 16'h736c, 16'h736c, 16'h734c, 16'h6b2c, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h6b4c, 16'h6b4c, 16'h736c, 16'h734c, 16'h734c, 16'h734c, 16'h736c, 16'h736c, 16'h734d, 16'h734c, 16'h732c, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h736c, 16'h7b8d, 16'h7b6d, 16'h7b6d, 16'h7b8d, 16'h736c, 16'h734c, 16'h6bc, 16'h63c, 16'h63c, 16'h63c, 16'h6b2c, 16'h6b2c, 16'h6b2c, 16'h6b4c, 16'h736c, 16'h736c, 16'h736d, 16'h736c, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h732c, 16'h734c, 16'h7b6c, 16'h942f, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc553, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha46f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9ce, 16'h9ce, 16'h7b2b, 16'h3944, 16'h20c2, 16'h20c2, 16'h20c2, 16'h20c2, 16'h1081, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'ha4b2, 16'ha4b3, 16'had14, 16'had14, 16'had14, 16'hb555, 16'hbd75, 16'hbd55, 16'hb514, 16'hb554, 16'hc595, 16'hc595, 16'hbd55, 16'hb534, 16'hbd54, 16'hb533, 16'had13, 16'hb574, 16'hbd74, 16'hbd95, 16'had12, 16'h7bad, 16'h732c, 16'h6aeb, 16'h62ea, 16'h734c, 16'hb553, 16'h83cd, 16'h2944, 16'h10a2, 16'h840, 16'h840, 16'h840, 16'h840, 16'h840, 16'h840, 16'h840, 16'h840, 16'h840, 16'h840, 16'h840, 16'h040, 16'h840, 16'h840, 16'h040, 16'h040, 16'h040, 16'h840, 16'h840, 16'h840, 16'h040, 16'h040, 16'h040, 16'h841, 16'h1081, 16'h4a48, 16'h62ca, 16'h6bb, 16'h62eb, 16'h528a, 16'h528a, 16'h6bc, 16'h736d, 16'h7b6d, 16'h736c, 16'h736c, 16'h736c, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h6b4c, 16'h734c, 16'h736c, 16'h736c, 16'h734c, 16'h736c, 16'h736c, 16'h7b6d, 16'h736d, 16'h734c, 16'h732c, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h736d, 16'h7b6d, 16'h7b8d, 16'h7b6d, 16'h7b6d, 16'h736c, 16'h734c, 16'h734c, 16'h734c, 16'h736c, 16'h734c, 16'h736c, 16'h734c, 16'h734c, 16'h736c, 16'h736c, 16'h736d, 16'h736d, 16'h736d, 16'h736d, 16'h736d, 16'h734c, 16'h734c, 16'h7b6c, 16'h7b6d, 16'h942f, 16'hc553, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc553, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd52, 16'hbd52, 16'hbd52, 16'hbd52, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hbd12, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9ce, 16'h9ce, 16'h7b2b, 16'h3144, 16'h20c2, 16'h20c2, 16'h20c2, 16'h20c2, 16'h1081, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h9c92, 16'ha4b2, 16'hacf3, 16'hacf3, 16'hb514, 16'hb555, 16'hb534, 16'hb514, 16'hb514, 16'hb554, 16'hbd55, 16'hc595, 16'hc5b6, 16'hc5b6, 16'hb554, 16'had13, 16'hb554, 16'hbd75, 16'hbd75, 16'hc5b5, 16'had12, 16'h7b8d, 16'h732c, 16'h6aeb, 16'h62eb, 16'h736d, 16'hb553, 16'h83cd, 16'h2944, 16'h10c2, 16'h841, 16'h841, 16'h840, 16'h840, 16'h840, 16'h840, 16'h840, 16'h840, 16'h840, 16'h840, 16'h840, 16'h040, 16'h840, 16'h040, 16'h040, 16'h040, 16'h040, 16'h840, 16'h840, 16'h840, 16'h840, 16'h040, 16'h841, 16'h841, 16'h1082, 16'h4a48, 16'h62ca, 16'h6bb, 16'h62eb, 16'h528a, 16'h528a, 16'h6bc, 16'h736d, 16'h736d, 16'h736c, 16'h736d, 16'h736d, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h6b4c, 16'h734c, 16'h736c, 16'h736c, 16'h734c, 16'h734c, 16'h736d, 16'h736d, 16'h736d, 16'h734c, 16'h732c, 16'h6b2c, 16'h6b4c, 16'h6b2c, 16'h6b2c, 16'h6b2c, 16'h736d, 16'h7bad, 16'h83cd, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h736c, 16'h734c, 16'h736c, 16'h736c, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h736d, 16'h736c, 16'h736d, 16'h736d, 16'h736d, 16'h736d, 16'h736c, 16'h734c, 16'h734c, 16'h7b6c, 16'h7b6d, 16'h942f, 16'hc553, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc553, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd52, 16'hbd52, 16'hbd52, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hacb0, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h94e, 16'h7b2b, 16'h3143, 16'h20e2, 16'h20c2, 16'h20c2, 16'h20c2, 16'h1081, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h9c91, 16'ha4b2, 16'ha4d3, 16'hacf3, 16'had14, 16'hb534, 16'hb555, 16'hb555, 16'hb534, 16'hb555, 16'hb554, 16'hbd75, 16'hbd95, 16'hc5d6, 16'hce17, 16'hc5b5, 16'hb533, 16'hbd75, 16'hbd95, 16'hc5d6, 16'hb532, 16'h7b8d, 16'h732c, 16'h6aeb, 16'h62eb, 16'h7b6d, 16'hb553, 16'h83cd, 16'h2923, 16'h10a2, 16'h840, 16'h841, 16'h840, 16'h840, 16'h840, 16'h840, 16'h040, 16'h840, 16'h840, 16'h840, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h840, 16'h840, 16'h840, 16'h841, 16'h840, 16'h840, 16'h841, 16'h1081, 16'h4a48, 16'h62ca, 16'h6bb, 16'h62eb, 16'h528a, 16'h528a, 16'h6bc, 16'h736c, 16'h736c, 16'h736c, 16'h736d, 16'h736d, 16'h734c, 16'h734c, 16'h734c, 16'h732c, 16'h6b2c, 16'h6b2c, 16'h734c, 16'h736c, 16'h736d, 16'h736c, 16'h734c, 16'h7b6d, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h734d, 16'h63c, 16'h63c, 16'h63c, 16'h6bc, 16'h6bc, 16'h7b6d, 16'h83cd, 16'h83ee, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h734c, 16'h734c, 16'h736c, 16'h736c, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h736d, 16'h736d, 16'h736d, 16'h736d, 16'h736d, 16'h736c, 16'h736d, 16'h736c, 16'h734c, 16'h7b6c, 16'h7b6d, 16'h942f, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd52, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h94e, 16'h7b2b, 16'h3143, 16'h20e2, 16'h20c2, 16'h20c2, 16'h20c2, 16'h1081, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h9471, 16'h9c92, 16'ha4b2, 16'ha4d3, 16'had13, 16'had14, 16'hb554, 16'hbd75, 16'hbd75, 16'hbd55, 16'hb555, 16'hbd75, 16'hbd75, 16'hbd95, 16'hcdf6, 16'hbd95, 16'hb533, 16'hbd95, 16'hc5b5, 16'hc5d6, 16'hb553, 16'h7b8d, 16'h734c, 16'h6bb, 16'h6bb, 16'h7b8d, 16'hb574, 16'h7bad, 16'h213, 16'h10a2, 16'h214, 16'h214, 16'h18e3, 16'h1881, 16'h1881, 16'h1081, 16'h841, 16'h840, 16'h840, 16'h840, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h840, 16'h840, 16'h841, 16'h1081, 16'h4a28, 16'h62cb, 16'h6aeb, 16'h62eb, 16'h528a, 16'h528a, 16'h6bc, 16'h736d, 16'h736c, 16'h736c, 16'h736c, 16'h736c, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h736c, 16'h736c, 16'h736c, 16'h736d, 16'h736d, 16'h7b8d, 16'h7bae, 16'h7bad, 16'h7bad, 16'h734d, 16'h63c, 16'h63c, 16'h63c, 16'h63c, 16'h6bc, 16'h7b8d, 16'h83cd, 16'h83ed, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h734c, 16'h734c, 16'h736c, 16'h736c, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h736d, 16'h736d, 16'h7b8d, 16'h736d, 16'h736d, 16'h736d, 16'h736d, 16'h736c, 16'h734c, 16'h7b6c, 16'h7b4c, 16'h942f, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc553, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hacd1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9c2f, 16'h9cf, 16'h9ce, 16'h7b2b, 16'h3144, 16'h20e2, 16'h20e2, 16'h20c2, 16'h20c2, 16'h1081, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h9430, 16'h9471, 16'h9c92, 16'ha4d2, 16'hacf3, 16'had13, 16'hb534, 16'hb554, 16'hbd75, 16'hc596, 16'hbd75, 16'hb555, 16'hbd55, 16'hbd95, 16'hbd75, 16'hbd74, 16'hc5b5, 16'hc5d6, 16'hc5b6, 16'hcdf6, 16'hbd94, 16'h83ad, 16'h7b8d, 16'h736d, 16'h734d, 16'h83ce, 16'hb574, 16'h7bac, 16'h20e3, 16'h3145, 16'h736d, 16'h738e, 16'h6b2b, 16'h6a66, 16'h626, 16'h3965, 16'h841, 16'h841, 16'h840, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h840, 16'h040, 16'h040, 16'h840, 16'h840, 16'h840, 16'h841, 16'h1081, 16'h4a48, 16'h62cb, 16'h6aeb, 16'h62eb, 16'h528a, 16'h528a, 16'h6bc, 16'h734c, 16'h736c, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h736c, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h736c, 16'h736c, 16'h736d, 16'h7b6d, 16'h7bad, 16'h83ad, 16'h83ae, 16'h7bae, 16'h736d, 16'h63c, 16'h63c, 16'h63c, 16'h6bc, 16'h6bc, 16'h7b8d, 16'h83cd, 16'h83ee, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h736c, 16'h734c, 16'h736c, 16'h736c, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h736d, 16'h736d, 16'h7b8d, 16'h736d, 16'h736d, 16'h736d, 16'h736d, 16'h736c, 16'h734c, 16'h736c, 16'h7b6d, 16'h9c2f, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc553, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha46f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9ce, 16'h94e, 16'h7b2b, 16'h3144, 16'h20e2, 16'h20c2, 16'h20c2, 16'h20c2, 16'h1081, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h8c2f, 16'h9450, 16'h9c71, 16'h9cb2, 16'ha4d2, 16'hacf3, 16'had14, 16'hb554, 16'hbd75, 16'hc595, 16'hc5b6, 16'hc5b6, 16'hbd75, 16'hbd95, 16'hc5b5, 16'hc5d6, 16'hcdd6, 16'hc5d6, 16'hc5d6, 16'hcdf6, 16'hc5b4, 16'ha4b1, 16'ha4b1, 16'ha4b1, 16'ha4b1, 16'ha4d1, 16'hb553, 16'h7bad, 16'h2924, 16'h3166, 16'h7b8e, 16'h7b8e, 16'h7b8e, 16'h734c, 16'h73c, 16'h39a7, 16'h841, 16'h841, 16'h840, 16'h840, 16'h840, 16'h840, 16'h040, 16'h040, 16'h040, 16'h040, 16'h041, 16'h040, 16'h040, 16'h040, 16'h840, 16'h840, 16'h840, 16'h841, 16'h1082, 16'h4a48, 16'h5aca, 16'h62eb, 16'h62cb, 16'h528a, 16'h528a, 16'h62eb, 16'h6b2c, 16'h6b2b, 16'h6b2c, 16'h734c, 16'h736c, 16'h736d, 16'h736d, 16'h736d, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h736c, 16'h736c, 16'h736d, 16'h7b6d, 16'h7bad, 16'h83ad, 16'h83ce, 16'h83ce, 16'h736d, 16'h63c, 16'h63c, 16'h63c, 16'h6bc, 16'h6b2c, 16'h7b8d, 16'h83cd, 16'h8bee, 16'h7b8d, 16'h7bad, 16'h7b8d, 16'h734c, 16'h734c, 16'h736c, 16'h736c, 16'h734c, 16'h734c, 16'h732c, 16'h734c, 16'h736d, 16'h736d, 16'h7b8d, 16'h736d, 16'h736d, 16'h736d, 16'h736d, 16'h736c, 16'h734c, 16'h736d, 16'h7b6d, 16'h942f, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha470, 16'ha470, 16'ha470, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9cf, 16'h94e, 16'h7b2b, 16'h3144, 16'h20e2, 16'h20c1, 16'h20c2, 16'h20c2, 16'h1081, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h83ef, 16'h8cf, 16'h9450, 16'h9c71, 16'h9cb2, 16'ha4d2, 16'hacf3, 16'had14, 16'hb534, 16'hb555, 16'hbd75, 16'hbd75, 16'hbd75, 16'hbd95, 16'hc5b6, 16'hc5b5, 16'hc5b5, 16'hc5b5, 16'hbd95, 16'hbd95, 16'hbd74, 16'hb553, 16'had33, 16'ha4d2, 16'h9cb1, 16'h9c70, 16'h944f, 16'h736c, 16'h41e7, 16'h3986, 16'h6b4d, 16'h6b4d, 16'h734d, 16'h734d, 16'h6b2d, 16'h39a6, 16'h1061, 16'h861, 16'h861, 16'h861, 16'h861, 16'h841, 16'h840, 16'h861, 16'h841, 16'h840, 16'h841, 16'h841, 16'h840, 16'h840, 16'h840, 16'h840, 16'h840, 16'h841, 16'h1082, 16'h4a48, 16'h62ca, 16'h6aeb, 16'h62eb, 16'h528a, 16'h528a, 16'h62eb, 16'h6b2b, 16'h6bb, 16'h6b2c, 16'h734c, 16'h736c, 16'h736d, 16'h736d, 16'h736c, 16'h7b8d, 16'h7bad, 16'h7bad, 16'h7b8d, 16'h736d, 16'h736d, 16'h7b6d, 16'h7b8d, 16'h7bad, 16'h83ae, 16'h83ce, 16'h83ce, 16'h736d, 16'h63c, 16'h63c, 16'h6bc, 16'h63c, 16'h6b2c, 16'h7b8d, 16'h83ce, 16'h8bee, 16'h838d, 16'h838d, 16'h7b8d, 16'h734c, 16'h734c, 16'h736c, 16'h736c, 16'h734c, 16'h734c, 16'h6b2c, 16'h734c, 16'h736d, 16'h736d, 16'h736d, 16'h736d, 16'h736d, 16'h736d, 16'h736d, 16'h734c, 16'h734c, 16'h734c, 16'h7b6c, 16'h942f, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc553, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd53, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hbd12, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h94e, 16'h7b4b, 16'h3144, 16'h20e2, 16'h20c2, 16'h20c2, 16'h20c2, 16'h1081, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h83ae, 16'h83ef, 16'h8c30, 16'h9451, 16'h9c71, 16'h9cb2, 16'ha4d2, 16'hacf3, 16'had13, 16'hb534, 16'hb554, 16'hb554, 16'hb554, 16'hbd55, 16'hbd75, 16'hbd75, 16'hbd75, 16'hb554, 16'hb554, 16'hb554, 16'hb554, 16'hb554, 16'had13, 16'ha4d2, 16'h9c70, 16'h942f, 16'h8bee, 16'h7bad, 16'h736c, 16'h6bb, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h6b2c, 16'h62ea, 16'h5a89, 16'h5a89, 16'h5a89, 16'h5a89, 16'h5289, 16'h4a28, 16'h426, 16'h4a6, 16'h3165, 16'h213, 16'h20e3, 16'h20e3, 16'h3164, 16'h3184, 16'h18c2, 16'h18c2, 16'h20e2, 16'h2124, 16'h3165, 16'h5a89, 16'h62ca, 16'h6aeb, 16'h62eb, 16'h528a, 16'h528a, 16'h62eb, 16'h6b2b, 16'h6bb, 16'h734c, 16'h734c, 16'h736d, 16'h736d, 16'h736c, 16'h736c, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h736c, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h7bae, 16'h83ae, 16'h83ae, 16'h736d, 16'h63c, 16'h63c, 16'h6bc, 16'h63c, 16'h6b2c, 16'h7b8d, 16'h83ad, 16'h8bee, 16'h838d, 16'h838d, 16'h7b8d, 16'h734c, 16'h734c, 16'h736c, 16'h736c, 16'h734c, 16'h6b4c, 16'h6b2b, 16'h6b2c, 16'h736d, 16'h736d, 16'h736d, 16'h736d, 16'h736d, 16'h736d, 16'h736d, 16'h734c, 16'h734c, 16'h734c, 16'h7b6d, 16'h942f, 16'hbd73, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc553, 16'hc553, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hbd12, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h94e, 16'h7b2a, 16'h3143, 16'h20e2, 16'h20c2, 16'h20c2, 16'h20c2, 16'h1081, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h83ef, 16'h8c10, 16'h9450, 16'h9c71, 16'h9cb2, 16'ha4d2, 16'ha4f3, 16'had13, 16'hb534, 16'hb554, 16'hb554, 16'hbd54, 16'hbd75, 16'hbd75, 16'hbd75, 16'hbd75, 16'hbd75, 16'hbd75, 16'hbd74, 16'hbd74, 16'hb554, 16'hb554, 16'hb554, 16'had33, 16'ha4d2, 16'h9c91, 16'h9450, 16'h8c2f, 16'h8ce, 16'h83ee, 16'h83cd, 16'h83ad, 16'h7bad, 16'h7bad, 16'h7bad, 16'h7bad, 16'h7bad, 16'h7bad, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h83ad, 16'h83ad, 16'h734c, 16'h736c, 16'h6ba, 16'h5aa9, 16'h62ea, 16'h5a88, 16'h3144, 16'h2923, 16'h3144, 16'h3985, 16'h41e7, 16'h5aaa, 16'h62aa, 16'h6aeb, 16'h62eb, 16'h528a, 16'h528a, 16'h62eb, 16'h6b2b, 16'h6b2b, 16'h6b2c, 16'h734c, 16'h736c, 16'h736d, 16'h736d, 16'h736d, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h7b6d, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h7bad, 16'h83ae, 16'h83ae, 16'h83ae, 16'h736d, 16'h62ec, 16'h63c, 16'h63c, 16'h63c, 16'h6b2c, 16'h7b8d, 16'h83cd, 16'h8bee, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h734c, 16'h734c, 16'h736c, 16'h736c, 16'h734c, 16'h6b4c, 16'h6b2c, 16'h6b2c, 16'h736d, 16'h736d, 16'h736d, 16'h736d, 16'h736d, 16'h736d, 16'h736d, 16'h736d, 16'h736c, 16'h736c, 16'h7b6c, 16'h942f, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc553, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha450, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h94e, 16'h7b2b, 16'h3143, 16'h20e2, 16'h20c2, 16'h20c2, 16'h20c2, 16'h1081, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h8c30, 16'h9450, 16'h9c91, 16'h9cb2, 16'ha4d2, 16'hacf3, 16'had13, 16'hb534, 16'hb554, 16'hb555, 16'hbd75, 16'hbd75, 16'hbd95, 16'hbd95, 16'hbd95, 16'hc595, 16'hbd95, 16'hbd95, 16'hbd95, 16'hbd95, 16'hbd75, 16'hbd74, 16'hb554, 16'hb554, 16'hb533, 16'ha4f2, 16'h9cb1, 16'h9450, 16'h8ce, 16'h83ee, 16'h83ee, 16'h83cd, 16'h83cd, 16'h7bad, 16'h7bad, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h7b8c, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h7b8c, 16'h736c, 16'h734b, 16'h62a9, 16'h3144, 16'h3123, 16'h3164, 16'h41c6, 16'h4a28, 16'h5aaa, 16'h5aaa, 16'h6aeb, 16'h62eb, 16'h528a, 16'h528a, 16'h62eb, 16'h6b2b, 16'h6b2c, 16'h734c, 16'h734c, 16'h736c, 16'h736d, 16'h736d, 16'h736c, 16'h7b8d, 16'h7b8d, 16'h738d, 16'h7b8d, 16'h736c, 16'h7b8c, 16'h7b8d, 16'h7b8d, 16'h7bad, 16'h83ae, 16'h83ce, 16'h83ce, 16'h736d, 16'h62ec, 16'h63c, 16'h63c, 16'h6bc, 16'h6b2c, 16'h7b8d, 16'h83ce, 16'h8bee, 16'h7b8d, 16'h7bad, 16'h7b8d, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h6b4c, 16'h6b2c, 16'h734c, 16'h736d, 16'h736d, 16'h736d, 16'h736d, 16'h736d, 16'h736d, 16'h736d, 16'h736d, 16'h734c, 16'h736c, 16'h7b6c, 16'h942f, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc553, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h94e, 16'h7b2b, 16'h3143, 16'h20e2, 16'h20e2, 16'h20c2, 16'h20c2, 16'h1081, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h9450, 16'h9471, 16'h9c92, 16'ha4b2, 16'ha4b2, 16'h9cb2, 16'ha4d3, 16'had13, 16'hb534, 16'hb554, 16'hb554, 16'hb574, 16'hb575, 16'hbd75, 16'hbd75, 16'hbd75, 16'hbd75, 16'hbd75, 16'hbd75, 16'hb554, 16'hb554, 16'hb554, 16'hb554, 16'had33, 16'ha4d2, 16'ha4b2, 16'h9cb1, 16'ha4b2, 16'h9450, 16'h8cf, 16'h83ce, 16'h83ce, 16'h83ce, 16'h83cd, 16'h83ad, 16'h7b8d, 16'h7b8d, 16'h7b6c, 16'h734c, 16'h732c, 16'h734b, 16'h734c, 16'h7b4c, 16'h7b6c, 16'h7b6c, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h62a9, 16'h3164, 16'h3143, 16'h39a5, 16'h5268, 16'h5248, 16'h5aaa, 16'h62aa, 16'h6bb, 16'h62eb, 16'h528a, 16'h528a, 16'h63b, 16'h734c, 16'h732c, 16'h734c, 16'h734c, 16'h736c, 16'h736c, 16'h736c, 16'h736c, 16'h736d, 16'h738d, 16'h734c, 16'h736c, 16'h7b6c, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h83ad, 16'h83ae, 16'h83ce, 16'h83cd, 16'h736d, 16'h63c, 16'h63c, 16'h6bc, 16'h6b2c, 16'h6b2c, 16'h7b8d, 16'h83ce, 16'h8bee, 16'h83ad, 16'h838d, 16'h7b8d, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h6b4c, 16'h734c, 16'h736c, 16'h736d, 16'h736d, 16'h736d, 16'h736d, 16'h736d, 16'h736c, 16'h734c, 16'h734c, 16'h736c, 16'h7b4c, 16'h942f, 16'hc553, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc553, 16'hc553, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hbd12, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hacd1, 16'hacd1, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb0, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha46f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9ce, 16'h7b2a, 16'h3143, 16'h20e2, 16'h20c2, 16'h20c2, 16'h20c2, 16'h1081, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h9c71, 16'h9c91, 16'h8cf, 16'h83ce, 16'h736d, 16'h83ce, 16'h9450, 16'h9c91, 16'h9cb2, 16'ha4b2, 16'ha4d2, 16'ha4f2, 16'hacf2, 16'hacf3, 16'hacf2, 16'ha4f2, 16'ha4f2, 16'ha4f2, 16'ha4f2, 16'ha4f2, 16'ha4f2, 16'ha4f2, 16'ha4d2, 16'h9c91, 16'h9471, 16'h9c91, 16'h9450, 16'h9c91, 16'h9c71, 16'h9450, 16'h8cf, 16'h83ad, 16'h7b8d, 16'h736c, 16'h732b, 16'h6bb, 16'h6bb, 16'h6aea, 16'h62ca, 16'h6aca, 16'h6aea, 16'h6aea, 16'h6aca, 16'h5a48, 16'h5a89, 16'h6aea, 16'h6bb, 16'h732b, 16'h736c, 16'h62ca, 16'h3964, 16'h3164, 16'h41c6, 16'h5a89, 16'h5249, 16'h62aa, 16'h62ca, 16'h6aeb, 16'h62eb, 16'h528a, 16'h528a, 16'h6bb, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h736c, 16'h736c, 16'h736c, 16'h736d, 16'h738d, 16'h734c, 16'h736d, 16'h736c, 16'h7b6d, 16'h7b8d, 16'h7b8d, 16'h83ad, 16'h83ce, 16'h83ce, 16'h83ae, 16'h736d, 16'h62ec, 16'h63c, 16'h6bc, 16'h6b2c, 16'h6b2c, 16'h7b8d, 16'h83cd, 16'h8bee, 16'h83ad, 16'h7bad, 16'h7b8d, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h6b2c, 16'h6b4c, 16'h734c, 16'h734d, 16'h734d, 16'h734d, 16'h734d, 16'h736d, 16'h736c, 16'h736c, 16'h734d, 16'h736c, 16'h7b4d, 16'h94f, 16'hc553, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc553, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hbd12, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hacb0, 16'h73b, 16'h527, 16'h5a69, 16'h93ee, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c2e, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h94e, 16'h7b2b, 16'h3143, 16'h20e2, 16'h20c2, 16'h20c2, 16'h20c2, 16'h1081, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h9cb1, 16'h8c2f, 16'h39c6, 16'h3165, 16'h41c7, 16'h4a8, 16'h5249, 16'h5269, 16'h5269, 16'h5269, 16'h5a89, 16'h5a8a, 16'h5a8a, 16'h5a89, 16'h5aaa, 16'h62ca, 16'h62ca, 16'h6bb, 16'h6b2c, 16'h6bb, 16'h62ca, 16'h62ca, 16'h62ca, 16'h62ca, 16'h5a8a, 16'h5a49, 16'h5a89, 16'h62ca, 16'h5a89, 16'h62ca, 16'h62aa, 16'h62a9, 16'h5a49, 16'h5a8, 16'h4165, 16'h3944, 16'h49c6, 16'h51e7, 16'h51e7, 16'h51e7, 16'h51c7, 16'h51e7, 16'h4985, 16'h394, 16'h5a48, 16'h6bb, 16'h732c, 16'h736c, 16'h7b8c, 16'h6bb, 16'h3985, 16'h3964, 16'h41e6, 16'h5a89, 16'h5269, 16'h62ca, 16'h62ca, 16'h6bb, 16'h62eb, 16'h528a, 16'h528a, 16'h6bb, 16'h734c, 16'h734c, 16'h6b2c, 16'h732c, 16'h732c, 16'h734c, 16'h734c, 16'h736c, 16'h736c, 16'h738d, 16'h736c, 16'h734c, 16'h736c, 16'h7b6d, 16'h7b8d, 16'h7b8d, 16'h83ae, 16'h83ce, 16'h83ce, 16'h83ae, 16'h736d, 16'h63c, 16'h63c, 16'h63c, 16'h6b2c, 16'h6b2c, 16'h7b8d, 16'h83cd, 16'h8bee, 16'h83ad, 16'h7bad, 16'h7b8d, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h6b4c, 16'h6b4c, 16'h6b2c, 16'h6b2c, 16'h734c, 16'h736c, 16'h734d, 16'h736d, 16'h734c, 16'h736d, 16'h736d, 16'h734c, 16'h734c, 16'h7b6d, 16'h7b6d, 16'h942f, 16'hc553, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc553, 16'hc553, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hacd1, 16'h62a9, 16'h293, 16'h20e3, 16'h20e3, 16'h49e7, 16'h94e, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h7b2a, 16'h3143, 16'h20e2, 16'h20e2, 16'h20c2, 16'h20c2, 16'h1081, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'ha4d2, 16'h8cf, 16'h2924, 16'h20e3, 16'h2945, 16'h39a6, 16'h4a8, 16'h5269, 16'h5269, 16'h4a28, 16'h4a28, 16'h4a48, 16'h5269, 16'h5269, 16'h5269, 16'h5269, 16'h5aa9, 16'h5a69, 16'h5249, 16'h5269, 16'h5228, 16'h527, 16'h51e7, 16'h49e7, 16'h49e7, 16'h4965, 16'h3944, 16'h3124, 16'h28e3, 16'h49c6, 16'h5a48, 16'h62aa, 16'h6aca, 16'h6aaa, 16'h5a48, 16'h49e7, 16'h6248, 16'h6269, 16'h6289, 16'h6aa9, 16'h6aa9, 16'h6aca, 16'h6269, 16'h51e7, 16'h6aaa, 16'h7b8d, 16'h83ad, 16'h83cd, 16'h83cd, 16'h734b, 16'h41a5, 16'h3984, 16'h41e6, 16'h5aa9, 16'h5269, 16'h62ca, 16'h62cb, 16'h6bb, 16'h62eb, 16'h528a, 16'h528a, 16'h62eb, 16'h734c, 16'h734b, 16'h6bb, 16'h6bb, 16'h6bb, 16'h6bb, 16'h6b2b, 16'h6b2b, 16'h6b4c, 16'h734c, 16'h6b4c, 16'h6b2b, 16'h734c, 16'h736c, 16'h7b8d, 16'h7b8d, 16'h83ad, 16'h83ce, 16'h83ae, 16'h83ae, 16'h736d, 16'h63c, 16'h63c, 16'h63c, 16'h6bc, 16'h6bc, 16'h736d, 16'h83cd, 16'h8bee, 16'h838d, 16'h7b8d, 16'h7b8d, 16'h734c, 16'h734c, 16'h734c, 16'h6b4c, 16'h6b4c, 16'h6b4c, 16'h6b2c, 16'h6b2c, 16'h6b4c, 16'h734c, 16'h734d, 16'h734d, 16'h734d, 16'h736d, 16'h736d, 16'h736c, 16'h734c, 16'h7b6c, 16'h7b6c, 16'h942f, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc574, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc553, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hb512, 16'hb512, 16'h836c, 16'h293, 16'h20e3, 16'h18e3, 16'h18e3, 16'h293, 16'h5a69, 16'hacb1, 16'hb4f1, 16'hb4f1, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hacb0, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha450, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h7b2a, 16'h3143, 16'h20e2, 16'h20c2, 16'h20c2, 16'h20c2, 16'h1081, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'hacf2, 16'h9c91, 16'h39a6, 16'h39c6, 16'h5acb, 16'h7b8d, 16'h8bef, 16'h9430, 16'h9430, 16'h8cf, 16'h8bef, 16'h8bef, 16'h942f, 16'h942f, 16'h942f, 16'h8bee, 16'h83ce, 16'h83ad, 16'h83ae, 16'h83ee, 16'h83ee, 16'h83ce, 16'h83ad, 16'h838d, 16'h838d, 16'h7b4c, 16'h6aaa, 16'h527, 16'h5228, 16'h6bb, 16'h83ad, 16'h836d, 16'h7bb, 16'h7b8d, 16'h7b8d, 16'h83ad, 16'h8bef, 16'h8bef, 16'h8bef, 16'h8bee, 16'h8bce, 16'h8bce, 16'h8bee, 16'h8bee, 16'h8bee, 16'h8bee, 16'h83ee, 16'h83ee, 16'h83ee, 16'h734b, 16'h41a5, 16'h3984, 16'h41e6, 16'h5a69, 16'h5269, 16'h62ca, 16'h62eb, 16'h6bb, 16'h62eb, 16'h528a, 16'h528a, 16'h62eb, 16'h734c, 16'h732b, 16'h6aea, 16'h62ea, 16'h6aea, 16'h6aeb, 16'h62eb, 16'h62eb, 16'h6bb, 16'h734c, 16'h734c, 16'h6bb, 16'h6b2c, 16'h734c, 16'h736c, 16'h7b8d, 16'h7bad, 16'h83ae, 16'h83ad, 16'h83ad, 16'h736d, 16'h63c, 16'h63c, 16'h63c, 16'h6bc, 16'h6b2c, 16'h736d, 16'h83ad, 16'h8bee, 16'h7bad, 16'h7b8d, 16'h7b8d, 16'h734c, 16'h734c, 16'h734c, 16'h6b4c, 16'h6b4c, 16'h6b4c, 16'h6b4c, 16'h6b2c, 16'h6b4c, 16'h6b4c, 16'h734d, 16'h734d, 16'h734d, 16'h734d, 16'h734c, 16'h734c, 16'h734c, 16'h7b6d, 16'h7b6d, 16'h94f, 16'hc573, 16'hc574, 16'hc574, 16'hc574, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc553, 16'hc553, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hb512, 16'hacd1, 16'h5227, 16'h20e3, 16'h18c2, 16'h18c2, 16'h18e3, 16'h20e3, 16'h294, 16'h8bcd, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha450, 16'ha450, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9ce, 16'h7b2b, 16'h3143, 16'h20c2, 16'h20c2, 16'h20c2, 16'h20c2, 16'h1061, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'had13, 16'hacf2, 16'h83ae, 16'h83ef, 16'h9cb1, 16'ha4d2, 16'ha4f2, 16'ha4f2, 16'ha4d2, 16'ha4d2, 16'ha4b2, 16'ha4b2, 16'ha4b2, 16'h9cb1, 16'h9c91, 16'h9c71, 16'h9c71, 16'h9c71, 16'h9c70, 16'h9c70, 16'h9c71, 16'h9c71, 16'h9450, 16'h9450, 16'h9450, 16'h9450, 16'h94f, 16'h83ad, 16'h8bee, 16'h942f, 16'h9470, 16'h9c70, 16'h94f, 16'h9c70, 16'h9c91, 16'h9c91, 16'h9c71, 16'h9c70, 16'h9470, 16'h9450, 16'h9450, 16'h9450, 16'h9450, 16'h9430, 16'h942f, 16'h942f, 16'h8c2f, 16'h8cf, 16'h8ce, 16'h736c, 16'h41c6, 16'h3984, 16'h41e6, 16'h4a28, 16'h5248, 16'h62ca, 16'h6aeb, 16'h6bc, 16'h62eb, 16'h526a, 16'h528a, 16'h62eb, 16'h734c, 16'h6b2b, 16'h62ea, 16'h62ca, 16'h6aea, 16'h62ea, 16'h5aaa, 16'h5aaa, 16'h6bb, 16'h734c, 16'h734c, 16'h6b2b, 16'h6b2c, 16'h736c, 16'h736c, 16'h7b6d, 16'h7bad, 16'h83ad, 16'h83ad, 16'h83ad, 16'h736d, 16'h63c, 16'h63c, 16'h63c, 16'h63c, 16'h6b2c, 16'h736d, 16'h83ad, 16'h8bee, 16'h7b8d, 16'h7b8d, 16'h7b8d, 16'h6b4c, 16'h6b2c, 16'h734c, 16'h6b4c, 16'h6b2c, 16'h6b4c, 16'h6b2c, 16'h6b2c, 16'h6b2c, 16'h6b2c, 16'h6b4c, 16'h6b4c, 16'h6b4c, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h7b6c, 16'h7b6d, 16'h942f, 16'hc573, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc553, 16'hc573, 16'hc553, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hb512, 16'h9c4f, 16'h3964, 16'h18e3, 16'h18e3, 16'h20e3, 16'h213, 16'h213, 16'h20e3, 16'h6aca, 16'hb4d1, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha450, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h94e, 16'h7b2a, 16'h3143, 16'h20c2, 16'h20c2, 16'h20c2, 16'h20c2, 16'h1061, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'hb553, 16'hb554, 16'hb554, 16'hb554, 16'hb534, 16'hb533, 16'had33, 16'had33, 16'had13, 16'had13, 16'had13, 16'had13, 16'hacf2, 16'ha4f2, 16'ha4f2, 16'ha4f2, 16'ha4f2, 16'ha4f2, 16'ha4f2, 16'ha4d2, 16'ha4f2, 16'ha4d2, 16'ha4d2, 16'ha4d1, 16'ha4d2, 16'ha4d2, 16'ha4d2, 16'ha4d2, 16'ha4b2, 16'ha4b1, 16'ha4b1, 16'ha4b2, 16'ha4b2, 16'ha4b1, 16'ha4b1, 16'ha4b2, 16'ha4b2, 16'ha4b1, 16'h9cb1, 16'h9c91, 16'h9c91, 16'h9c70, 16'h9c70, 16'h9450, 16'h9450, 16'h9450, 16'h9450, 16'h944f, 16'h942f, 16'h7b8d, 16'h41c6, 16'h39a5, 16'h4a6, 16'h4a28, 16'h5248, 16'h62aa, 16'h62ca, 16'h62ca, 16'h5aaa, 16'h4a29, 16'h4a29, 16'h5289, 16'h62ca, 16'h5aa9, 16'h5248, 16'h5248, 16'h5248, 16'h5248, 16'h5269, 16'h5a89, 16'h62cb, 16'h6b2c, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h736c, 16'h736d, 16'h7bad, 16'h83ae, 16'h83ae, 16'h83ad, 16'h736d, 16'h63b, 16'h63c, 16'h63c, 16'h63c, 16'h6b2c, 16'h736c, 16'h83ad, 16'h8bee, 16'h7b8d, 16'h7b8d, 16'h7b6d, 16'h6b2c, 16'h6b2b, 16'h6b2c, 16'h6b4c, 16'h6b2c, 16'h6b2c, 16'h6b2c, 16'h6b2c, 16'h6b2c, 16'h6b2c, 16'h6b2c, 16'h6b2c, 16'h6b4c, 16'h736c, 16'h734c, 16'h734c, 16'h734c, 16'h7b6d, 16'h7b6d, 16'h942f, 16'hc573, 16'hc594, 16'hc574, 16'hc574, 16'hc574, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc553, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hb512, 16'h8bed, 16'h2924, 16'h18e3, 16'h20e3, 16'h214, 16'h213, 16'h20e3, 16'h20e3, 16'h4a28, 16'hacd1, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb0, 16'hacb0, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9ce, 16'h7b2a, 16'h3143, 16'h20c1, 16'h20c2, 16'h20c2, 16'h20c2, 16'h1081, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'hb554, 16'hb554, 16'hb553, 16'hb533, 16'had13, 16'hacf2, 16'hacf2, 16'had13, 16'had13, 16'had13, 16'had13, 16'had12, 16'hacf2, 16'ha4f2, 16'ha4f2, 16'ha4d2, 16'ha4f2, 16'ha4f2, 16'ha4f2, 16'ha4f2, 16'ha4d2, 16'ha4d2, 16'ha4b2, 16'ha4d2, 16'ha4d2, 16'ha4d2, 16'ha4d2, 16'ha4f2, 16'ha4f2, 16'ha4f2, 16'ha4d2, 16'ha4d2, 16'ha4d2, 16'ha4d2, 16'ha4b2, 16'ha4d2, 16'ha4b2, 16'ha4b2, 16'h9cb1, 16'h9cb1, 16'h9c91, 16'h9470, 16'h83ae, 16'h6bb, 16'h62ea, 16'h5aaa, 16'h5289, 16'h5248, 16'h4a28, 16'h41c6, 16'h20e3, 16'h18c2, 16'h20e3, 16'h213, 16'h20e3, 16'h213, 16'h20e3, 16'h20e3, 16'h18e3, 16'h18c3, 16'h18c3, 16'h20e3, 16'h20e3, 16'h20e3, 16'h18e3, 16'h213, 16'h2944, 16'h2944, 16'h39a6, 16'h41e7, 16'h5289, 16'h6b2c, 16'h734c, 16'h734c, 16'h6b2c, 16'h734c, 16'h734c, 16'h736c, 16'h7b8d, 16'h7bad, 16'h7bad, 16'h7b8d, 16'h736d, 16'h62ec, 16'h63c, 16'h63c, 16'h63c, 16'h6bc, 16'h736c, 16'h83ad, 16'h83ce, 16'h7b6d, 16'h7b6d, 16'h736c, 16'h732c, 16'h6b2b, 16'h6b2b, 16'h6b2c, 16'h6b2c, 16'h6b2c, 16'h6b2c, 16'h6bc, 16'h63c, 16'h6b2c, 16'h6b2c, 16'h6b2c, 16'h6b2c, 16'h6b4c, 16'h734c, 16'h734c, 16'h734c, 16'h7b4c, 16'h7b6d, 16'h94f, 16'hc573, 16'hc594, 16'hc594, 16'hc594, 16'hc574, 16'hc574, 16'hc574, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc553, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'h838c, 16'h213, 16'h18e2, 16'h18e3, 16'h213, 16'h213, 16'h20e3, 16'h20e3, 16'h41c6, 16'hacb1, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h7b2a, 16'h3143, 16'h20c1, 16'h20c2, 16'h20c2, 16'h20c2, 16'h1081, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'hb554, 16'hb533, 16'h9c2e, 16'h834b, 16'h7b2a, 16'h838b, 16'h94d, 16'h9c4e, 16'h9c4e, 16'h9c4e, 16'h9c4f, 16'h9c4f, 16'h9c6f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c4f, 16'h9c4f, 16'h9c4e, 16'h93ed, 16'h83ac, 16'h83ce, 16'h942f, 16'h9c90, 16'h9c90, 16'h9cb1, 16'ha4d2, 16'ha4d2, 16'ha4f2, 16'ha4d2, 16'ha4d2, 16'ha4d2, 16'ha4d2, 16'ha4d2, 16'ha4d2, 16'ha4d2, 16'h9cb1, 16'h8cf, 16'h736c, 16'h62ca, 16'h5a89, 16'h5248, 16'h41c7, 16'h39a5, 16'h2964, 16'h18e3, 16'h1082, 16'h861, 16'h861, 16'h861, 16'h861, 16'h861, 16'h861, 16'h1082, 16'h10a2, 16'h18a2, 16'h18c2, 16'h18c3, 16'h18c3, 16'h18e3, 16'h20e3, 16'h213, 16'h213, 16'h214, 16'h213, 16'h20e3, 16'h20e3, 16'h18c2, 16'h18c2, 16'h18a2, 16'h3185, 16'h6bb, 16'h6b4c, 16'h6b4c, 16'h62eb, 16'h6bb, 16'h6bc, 16'h6bc, 16'h6b2c, 16'h6b2c, 16'h734c, 16'h734c, 16'h6b2c, 16'h62eb, 16'h62ec, 16'h62ec, 16'h63c, 16'h63c, 16'h734c, 16'h7b8d, 16'h7bad, 16'h7b6d, 16'h736d, 16'h736c, 16'h6b2c, 16'h6b2b, 16'h6b2b, 16'h6b2c, 16'h6b2c, 16'h6b2c, 16'h6b2c, 16'h6bc, 16'h62ec, 16'h62ec, 16'h6bc, 16'h6b2c, 16'h6b2c, 16'h6b2c, 16'h6b4c, 16'h6b2c, 16'h734c, 16'h7b6c, 16'h7b6c, 16'h942f, 16'hc573, 16'hc594, 16'hc594, 16'hc594, 16'hc594, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc573, 16'hc573, 16'hc553, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'h83ad, 16'h293, 16'h18c2, 16'h18c3, 16'h20e3, 16'h213, 16'h213, 16'h213, 16'h39a6, 16'ha490, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h732a, 16'h3143, 16'h20c2, 16'h20c2, 16'h20c2, 16'h20c2, 16'h1081, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'hb554, 16'hacf2, 16'h8b29, 16'h61c5, 16'h59c6, 16'h7268, 16'h82ea, 16'h8b2b, 16'h8b4b, 16'h8b6b, 16'h8b6b, 16'h832a, 16'h7ae9, 16'h7ba, 16'h832a, 16'h832a, 16'h832a, 16'h83a, 16'h7aa9, 16'h7268, 16'h6288, 16'h62ca, 16'h736c, 16'h8c2e, 16'h9470, 16'h9c91, 16'ha4b1, 16'ha4d2, 16'ha4d2, 16'ha4d2, 16'ha4d2, 16'ha4d2, 16'ha4d2, 16'ha4b2, 16'ha4b2, 16'h9c91, 16'h734c, 16'h4a28, 16'h39a6, 16'h3185, 16'h3185, 16'h3165, 16'h2944, 16'h3185, 16'h3185, 16'h18c2, 16'h1082, 16'h1082, 16'h2944, 16'h3185, 16'h214, 16'h18e3, 16'h10a2, 16'h1081, 16'h2944, 16'h3185, 16'h3186, 16'h3185, 16'h3165, 16'h2945, 16'h3185, 16'h39a6, 16'h41c7, 16'h41e7, 16'h41c6, 16'h39c6, 16'h39c6, 16'h41c6, 16'h41c6, 16'h39c6, 16'h4a28, 16'h6bb, 16'h734c, 16'h6b2c, 16'h62eb, 16'h63c, 16'h63c, 16'h63c, 16'h5acc, 16'h62eb, 16'h63b, 16'h6bb, 16'h62eb, 16'h5aab, 16'h52ab, 16'h52ab, 16'h5aab, 16'h5aab, 16'h62eb, 16'h63c, 16'h6bc, 16'h6b2c, 16'h6b2c, 16'h6b2c, 16'h6b2c, 16'h6b2c, 16'h6b2c, 16'h6b2c, 16'h6b2c, 16'h6b2c, 16'h6b2c, 16'h6bc, 16'h62ec, 16'h62ec, 16'h63c, 16'h63c, 16'h6b2c, 16'h6b2c, 16'h6b2c, 16'h6b2c, 16'h734c, 16'h734d, 16'h7b6d, 16'h942f, 16'hc574, 16'hc594, 16'hc594, 16'hc594, 16'hc594, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc573, 16'hc573, 16'hc573, 16'hc553, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'h8bcd, 16'h2924, 16'h18c3, 16'h18e3, 16'h213, 16'h214, 16'h214, 16'h213, 16'h4a7, 16'hacb1, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h732b, 16'h3123, 16'h20c2, 16'h20c2, 16'h20c2, 16'h20c2, 16'h1081, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'hb554, 16'ha4f2, 16'h5a27, 16'h30e3, 16'h30e3, 16'h4144, 16'h49c6, 16'h59e7, 16'h5a7, 16'h6248, 16'h6268, 16'h5a7, 16'h51a6, 16'h51e7, 16'h5a28, 16'h6247, 16'h6247, 16'h6247, 16'h6227, 16'h4965, 16'h3964, 16'h5248, 16'h6b2b, 16'h83ce, 16'h8c2f, 16'h9450, 16'h9c91, 16'h9cb1, 16'h9cb1, 16'h9c91, 16'h9c91, 16'h9c91, 16'h9c71, 16'h9470, 16'h9450, 16'h7b6d, 16'h4a7, 16'h39a6, 16'h3985, 16'h3185, 16'h3165, 16'h3164, 16'h2944, 16'h2124, 16'h213, 16'h18e2, 16'h18c2, 16'h10a2, 16'h4a48, 16'h6b2b, 16'h5248, 16'h41e6, 16'h2924, 16'h20e3, 16'h5289, 16'h62ea, 16'h5aca, 16'h5aa9, 16'h5248, 16'h4a28, 16'h5269, 16'h5aaa, 16'h6aeb, 16'h6bb, 16'h62ea, 16'h62ca, 16'h62aa, 16'h62aa, 16'h5a89, 16'h5269, 16'h5aaa, 16'h6b2c, 16'h734c, 16'h6b2c, 16'h62eb, 16'h63c, 16'h63c, 16'h62ec, 16'h5acb, 16'h62eb, 16'h63b, 16'h63b, 16'h62eb, 16'h52aa, 16'h52aa, 16'h528b, 16'h52aa, 16'h5aaa, 16'h5acb, 16'h62eb, 16'h62ec, 16'h63c, 16'h63c, 16'h6bc, 16'h6b2b, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h6b4c, 16'h6bc, 16'h6b2c, 16'h6b2c, 16'h63c, 16'h6bc, 16'h63b, 16'h63b, 16'h63b, 16'h6bc, 16'h734c, 16'h734c, 16'h942f, 16'hc574, 16'hc594, 16'hc594, 16'hc594, 16'hc594, 16'hc594, 16'hc594, 16'hc594, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc573, 16'hc573, 16'hc573, 16'hc553, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd32, 16'h9c4f, 16'h3164, 16'h20e3, 16'h20e3, 16'h213, 16'h213, 16'h213, 16'h2924, 16'h62a9, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c2e, 16'h7b2b, 16'h3143, 16'h20c2, 16'h20c2, 16'h20e2, 16'h20c2, 16'h1081, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'hb554, 16'ha4f2, 16'h4a28, 16'h20a2, 16'h18a2, 16'h213, 16'h3144, 16'h3985, 16'h39a6, 16'h41a6, 16'h3985, 16'h3144, 16'h3144, 16'h3965, 16'h39a5, 16'h49e6, 16'h5227, 16'h527, 16'h49e6, 16'h3124, 16'h2924, 16'h49e6, 16'h5248, 16'h62a9, 16'h6aca, 16'h73b, 16'h73b, 16'h6aeb, 16'h73b, 16'h732b, 16'h72eb, 16'h6aca, 16'h6289, 16'h5a48, 16'h5a69, 16'h5248, 16'h41c6, 16'h3986, 16'h3185, 16'h3165, 16'h3164, 16'h2944, 16'h2944, 16'h2124, 16'h2123, 16'h213, 16'h18e3, 16'h10a2, 16'h3985, 16'h62ea, 16'h5a89, 16'h4a27, 16'h3985, 16'h3185, 16'h5269, 16'h3185, 16'h213, 16'h2924, 16'h39c6, 16'h39c6, 16'h4a28, 16'h5aa9, 16'h6aea, 16'h6bb, 16'h6aea, 16'h62ca, 16'h62ca, 16'h62aa, 16'h5a89, 16'h5269, 16'h62ca, 16'h6b2c, 16'h734c, 16'h6b2c, 16'h62eb, 16'h62eb, 16'h63c, 16'h62ec, 16'h62eb, 16'h62eb, 16'h6bb, 16'h6bb, 16'h62cb, 16'h52aa, 16'h528a, 16'h528a, 16'h52aa, 16'h52aa, 16'h5acb, 16'h5aeb, 16'h62ec, 16'h63c, 16'h6bc, 16'h6bc, 16'h6b2c, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h736c, 16'h6b4c, 16'h6b2b, 16'h6b2b, 16'h6b2c, 16'h63b, 16'h6bc, 16'h63b, 16'h63b, 16'h62eb, 16'h6b2c, 16'h736d, 16'h7b6c, 16'h942f, 16'hc594, 16'hcd94, 16'hcd94, 16'hcd94, 16'hcd94, 16'hcd94, 16'hc594, 16'hc594, 16'hc594, 16'hc594, 16'hc574, 16'hc574, 16'hc574, 16'hc573, 16'hc573, 16'hc573, 16'hc553, 16'hc553, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd33, 16'hbd33, 16'hacd1, 16'h5227, 16'h213, 16'h20e3, 16'h18e3, 16'h18e3, 16'h213, 16'h4a28, 16'h8b8d, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h7b2b, 16'h3143, 16'h20c2, 16'h20c2, 16'h20e2, 16'h20c2, 16'h1061, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'hb554, 16'hacf2, 16'h72a9, 16'h38e3, 16'h3124, 16'h49c6, 16'h5a7, 16'h6248, 16'h5a28, 16'h6269, 16'h6269, 16'h5a28, 16'h5a28, 16'h527, 16'h5228, 16'h5a28, 16'h51e7, 16'h51e7, 16'h51e7, 16'h51c7, 16'h51c6, 16'h51c6, 16'h51c6, 16'h51c6, 16'h59e7, 16'h59e7, 16'h51c6, 16'h49c6, 16'h5a7, 16'h6aa9, 16'h6289, 16'h4185, 16'h3945, 16'h3944, 16'h41a6, 16'h4a7, 16'h39a6, 16'h3185, 16'h3165, 16'h3164, 16'h2944, 16'h2944, 16'h2924, 16'h2124, 16'h2123, 16'h213, 16'h20e3, 16'h18c2, 16'h18c2, 16'h4a27, 16'h5a89, 16'h4a28, 16'h3986, 16'h2944, 16'h31a5, 16'h10a2, 16'h1082, 16'h1081, 16'h18c2, 16'h18a2, 16'h2924, 16'h5269, 16'h6aeb, 16'h6bb, 16'h6aeb, 16'h62ca, 16'h62ca, 16'h62ca, 16'h5a89, 16'h5269, 16'h62ca, 16'h6b2c, 16'h6b4c, 16'h6b2b, 16'h62cb, 16'h5aeb, 16'h63c, 16'h63c, 16'h63c, 16'h63c, 16'h6bb, 16'h6bb, 16'h62cb, 16'h528a, 16'h528a, 16'h528a, 16'h528a, 16'h52aa, 16'h5aab, 16'h5aeb, 16'h62ec, 16'h63c, 16'h6bc, 16'h6b2c, 16'h6b2b, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h736c, 16'h734c, 16'h6b2c, 16'h6bc, 16'h6b2c, 16'h6b2c, 16'h6bc, 16'h6bb, 16'h63b, 16'h62eb, 16'h6b2c, 16'h7b6d, 16'h7b6c, 16'h942f, 16'hc594, 16'hcdb4, 16'hcd94, 16'hcd94, 16'hcd94, 16'hcd94, 16'hcd94, 16'hcd94, 16'hc594, 16'hc594, 16'hc594, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc573, 16'hc573, 16'hc573, 16'hc553, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd32, 16'h7b6c, 16'h2924, 16'h213, 16'h20e3, 16'h213, 16'h31a5, 16'h7b4c, 16'ha470, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'ha490, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h7b2b, 16'h3143, 16'h20c2, 16'h20c2, 16'h20e2, 16'h20c2, 16'h1081, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'hb554, 16'ha4b1, 16'h6a69, 16'h30c3, 16'h3124, 16'h49c7, 16'h5a69, 16'h62aa, 16'h62a9, 16'h62aa, 16'h62aa, 16'h6aaa, 16'h6acb, 16'h6aaa, 16'h628a, 16'h6289, 16'h5a48, 16'h5a48, 16'h5a48, 16'h5a48, 16'h6249, 16'h5a28, 16'h5a28, 16'h5a28, 16'h5a28, 16'h5a28, 16'h5a28, 16'h528, 16'h51e7, 16'h5a89, 16'h52ca, 16'h29a6, 16'h1944, 16'h2145, 16'h31a6, 16'h4a7, 16'h3986, 16'h3165, 16'h3144, 16'h3144, 16'h2944, 16'h2944, 16'h2924, 16'h2124, 16'h2123, 16'h213, 16'h20e3, 16'h18c2, 16'h1082, 16'h39a6, 16'h5a89, 16'h4a27, 16'h3985, 16'h2124, 16'h29c6, 16'h21c6, 16'h29c6, 16'h31a5, 16'h2944, 16'h18a2, 16'h213, 16'h5268, 16'h6aeb, 16'h62eb, 16'h6bb, 16'h62ea, 16'h62ca, 16'h62ca, 16'h5a89, 16'h5268, 16'h62ca, 16'h6b2c, 16'h6b2c, 16'h6b2c, 16'h5acb, 16'h5aec, 16'h62ec, 16'h63b, 16'h6b2c, 16'h6b2c, 16'h6bb, 16'h6bb, 16'h62cb, 16'h528a, 16'h528a, 16'h528a, 16'h528a, 16'h52aa, 16'h5acb, 16'h5aeb, 16'h62eb, 16'h63c, 16'h6bc, 16'h6b2c, 16'h6b2c, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h6b2c, 16'h6b2c, 16'h6b2c, 16'h6b2c, 16'h6b2c, 16'h63c, 16'h62eb, 16'h62eb, 16'h6bc, 16'h7b6d, 16'h7b6d, 16'h942f, 16'hc594, 16'hcdb4, 16'hcdb4, 16'hcdb4, 16'hcdb4, 16'hcdb4, 16'hcd94, 16'hcd94, 16'hcd94, 16'hc594, 16'hc594, 16'hc594, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc573, 16'hc573, 16'hc553, 16'hc553, 16'hc553, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'ha4b1, 16'h5248, 16'h2945, 16'h2924, 16'h2965, 16'h41c7, 16'h8bad, 16'hb4f2, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha450, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h7b2b, 16'h3143, 16'h20e2, 16'h20c2, 16'h20c2, 16'h20c2, 16'h1081, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'hb554, 16'hb513, 16'h8b2c, 16'h59a7, 16'h5a28, 16'h6aaa, 16'h7b2c, 16'h834d, 16'h834d, 16'h836d, 16'h836d, 16'h8b6d, 16'h8b4d, 16'h8b6d, 16'h936d, 16'h936d, 16'h8b6d, 16'h8b6d, 16'h8b6d, 16'h836d, 16'h8b8d, 16'h8b6d, 16'h836c, 16'h838d, 16'h8b8d, 16'h838d, 16'h8b8d, 16'h8b8d, 16'h7bb, 16'h4a28, 16'h3228, 16'h3a48, 16'h4269, 16'h4289, 16'h4aa9, 16'h427, 16'h3185, 16'h3165, 16'h3164, 16'h2944, 16'h2944, 16'h2944, 16'h2924, 16'h2924, 16'h2123, 16'h213, 16'h20e3, 16'h18c2, 16'h10a2, 16'h41e7, 16'h62a9, 16'h5248, 16'h3165, 16'h213, 16'h31e7, 16'h2a27, 16'h327, 16'h41e6, 16'h2944, 16'h213, 16'h39a6, 16'h5289, 16'h5aaa, 16'h5269, 16'h62ca, 16'h62ea, 16'h62ea, 16'h62ca, 16'h5a89, 16'h5268, 16'h62ca, 16'h6b4c, 16'h6b4c, 16'h6b2c, 16'h5acb, 16'h62ec, 16'h62eb, 16'h63c, 16'h6b2c, 16'h6b2c, 16'h6bb, 16'h6bb, 16'h62eb, 16'h528a, 16'h52aa, 16'h528a, 16'h528a, 16'h528a, 16'h5acb, 16'h62eb, 16'h62eb, 16'h63c, 16'h63c, 16'h6b2c, 16'h6b2c, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h6b2c, 16'h6bc, 16'h6bb, 16'h6bc, 16'h6bc, 16'h6bb, 16'h63b, 16'h62eb, 16'h62cb, 16'h6bb, 16'h7b6c, 16'h7b6d, 16'h942f, 16'hcdb4, 16'hcdb5, 16'hcdb5, 16'hcdb4, 16'hcdb4, 16'hcdb4, 16'hcdb4, 16'hcdb4, 16'hcd94, 16'hcd94, 16'hc594, 16'hc594, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc573, 16'hc573, 16'hc573, 16'hc553, 16'hc553, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'h942f, 16'h6aeb, 16'h5a69, 16'h41e7, 16'h62aa, 16'ha470, 16'hbd32, 16'hbd32, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha46f, 16'ha470, 16'ha470, 16'ha470, 16'ha450, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h7b2b, 16'h3123, 16'h20c2, 16'h20c2, 16'h20c2, 16'h20c2, 16'h1081, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'hb554, 16'hb554, 16'hacd2, 16'ha491, 16'ha4d2, 16'hacf2, 16'hacf3, 16'had13, 16'had13, 16'had13, 16'hacf3, 16'hacf2, 16'ha4d2, 16'ha4f2, 16'ha4d2, 16'ha4d2, 16'ha4d2, 16'ha4d2, 16'ha4b1, 16'ha4b1, 16'h9cb1, 16'h9c91, 16'h9c91, 16'h9c90, 16'h9c90, 16'h9c70, 16'h9c70, 16'h9c70, 16'h83ee, 16'h5269, 16'h3a28, 16'h5aeb, 16'h8c2f, 16'h944f, 16'h7bad, 16'h4a27, 16'h3185, 16'h3165, 16'h3164, 16'h3164, 16'h2944, 16'h2944, 16'h2924, 16'h2924, 16'h2923, 16'h213, 16'h20e3, 16'h18e2, 16'h18a2, 16'h5248, 16'h62aa, 16'h4a28, 16'h3164, 16'h20e3, 16'h4228, 16'h3248, 16'h3227, 16'h4a27, 16'h20e3, 16'h18a2, 16'h3185, 16'h5a89, 16'h5a89, 16'h5269, 16'h5aa9, 16'h62ea, 16'h62aa, 16'h5aaa, 16'h5269, 16'h5248, 16'h62ca, 16'h6b4c, 16'h6b2c, 16'h6b2b, 16'h5acb, 16'h62ec, 16'h62ec, 16'h63c, 16'h6b4c, 16'h6b2c, 16'h6b2b, 16'h6bb, 16'h62eb, 16'h52aa, 16'h52aa, 16'h52aa, 16'h528a, 16'h528a, 16'h5aaa, 16'h62eb, 16'h63c, 16'h6bc, 16'h6bc, 16'h6b2c, 16'h6b2c, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h6b2c, 16'h6bb, 16'h6bb, 16'h6bb, 16'h6bb, 16'h6bb, 16'h63b, 16'h63b, 16'h62eb, 16'h6bc, 16'h736c, 16'h7b6d, 16'h942f, 16'hcdb4, 16'hcdb5, 16'hcdb5, 16'hcdb5, 16'hcdb5, 16'hcdb5, 16'hcdb5, 16'hcdb4, 16'hcdb4, 16'hcd94, 16'hcd94, 16'hcd94, 16'hc594, 16'hc594, 16'hc594, 16'hc594, 16'hc574, 16'hc574, 16'hc574, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc553, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hacd1, 16'h94f, 16'h93ee, 16'hacd1, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h7b2b, 16'h3143, 16'h20e2, 16'h20e2, 16'h20c2, 16'h20c2, 16'h1081, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'hb554, 16'hb554, 16'hb554, 16'hb554, 16'hb554, 16'hb534, 16'hb534, 16'had33, 16'had33, 16'had13, 16'had13, 16'had13, 16'had13, 16'hacf2, 16'hacf2, 16'ha4f2, 16'ha4d2, 16'ha4d2, 16'ha4d2, 16'ha4d2, 16'ha4b2, 16'ha4b1, 16'h9cb1, 16'h9cb1, 16'h9c91, 16'h9c91, 16'h9c91, 16'h9c91, 16'h8ce, 16'h5a68, 16'h31e7, 16'h4248, 16'h62ea, 16'h942f, 16'h83ce, 16'h4a27, 16'h3185, 16'h3164, 16'h3164, 16'h3164, 16'h2944, 16'h2944, 16'h2944, 16'h2924, 16'h2923, 16'h213, 16'h213, 16'h18e2, 16'h18a2, 16'h5248, 16'h62aa, 16'h4a28, 16'h3144, 16'h18c2, 16'h3a27, 16'h3248, 16'h3227, 16'h427, 16'h18e2, 16'h1081, 16'h2964, 16'h5268, 16'h49e7, 16'h5aa9, 16'h5aa9, 16'h62ea, 16'h5aa9, 16'h5269, 16'h4a28, 16'h4a27, 16'h5aaa, 16'h6b4c, 16'h734c, 16'h6b2c, 16'h62cb, 16'h62eb, 16'h62eb, 16'h63b, 16'h734c, 16'h734c, 16'h6b2b, 16'h6bb, 16'h62ea, 16'h5aaa, 16'h52aa, 16'h52aa, 16'h52aa, 16'h528a, 16'h52aa, 16'h5acb, 16'h62eb, 16'h63c, 16'h6bc, 16'h6b2c, 16'h6b2c, 16'h734c, 16'h734c, 16'h736c, 16'h734c, 16'h734c, 16'h734c, 16'h6b2c, 16'h6bc, 16'h6bc, 16'h6bc, 16'h6bb, 16'h6bb, 16'h6bb, 16'h63b, 16'h62eb, 16'h6bb, 16'h734c, 16'h736c, 16'h9c2f, 16'hcdb5, 16'hcdd5, 16'hcdd5, 16'hcdd5, 16'hcdd5, 16'hcdd5, 16'hcdb5, 16'hcdb5, 16'hcdb4, 16'hcdb4, 16'hcdb4, 16'hcdb4, 16'hcd94, 16'hcd94, 16'hcd94, 16'hc594, 16'hc594, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc573, 16'hc573, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c2f, 16'h7b4b, 16'h3143, 16'h20e2, 16'h20e2, 16'h20c2, 16'h20c2, 16'h1081, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'hb554, 16'hb554, 16'hb534, 16'hb534, 16'had33, 16'had33, 16'had13, 16'had13, 16'hacf2, 16'hacf2, 16'ha4f2, 16'ha4d2, 16'ha4d2, 16'ha4d2, 16'ha4b1, 16'h9cb1, 16'h9c91, 16'ha4b2, 16'ha4d2, 16'ha4d2, 16'ha4d2, 16'ha4b2, 16'ha4b1, 16'h9cb1, 16'h9cb1, 16'h9cb1, 16'h9cb1, 16'h9c91, 16'h8ce, 16'h5268, 16'h39e7, 16'h52a9, 16'h41c6, 16'h62ca, 16'h83ee, 16'h4a27, 16'h3985, 16'h3164, 16'h3144, 16'h3144, 16'h3144, 16'h2944, 16'h2944, 16'h2924, 16'h2924, 16'h213, 16'h213, 16'h18e2, 16'h18a2, 16'h5248, 16'h62aa, 16'h4a27, 16'h2944, 16'h18c2, 16'h4227, 16'h3248, 16'h3227, 16'h427, 16'h18c2, 16'h861, 16'h2944, 16'h5269, 16'h5a89, 16'h62eb, 16'h5a89, 16'h62ea, 16'h5aaa, 16'h5248, 16'h427, 16'h41e7, 16'h5289, 16'h6b2b, 16'h6b4c, 16'h6b2c, 16'h62cb, 16'h62cb, 16'h5acb, 16'h62eb, 16'h6b4c, 16'h734c, 16'h6bb, 16'h6bb, 16'h62ea, 16'h52aa, 16'h52aa, 16'h52aa, 16'h52aa, 16'h528a, 16'h52aa, 16'h5acb, 16'h62eb, 16'h62ec, 16'h6bc, 16'h6b2c, 16'h6b2c, 16'h734c, 16'h734c, 16'h736c, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h6bb, 16'h6bc, 16'h6b2c, 16'h6bc, 16'h6bb, 16'h63b, 16'h63b, 16'h62eb, 16'h6b2b, 16'h736c, 16'h7b6c, 16'h9c30, 16'hcdd5, 16'hd5d5, 16'hd5d5, 16'hd5d5, 16'hd5d5, 16'hcdd5, 16'hcdd5, 16'hcdb5, 16'hcdb5, 16'hcdb5, 16'hcdb5, 16'hcdb5, 16'hcdb4, 16'hcdb4, 16'hcd94, 16'hcd94, 16'hcd94, 16'hcd94, 16'hc594, 16'hc594, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc553, 16'hc553, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h7b4b, 16'h3143, 16'h20e2, 16'h20e2, 16'h20c2, 16'h20c2, 16'h1081, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'ha4d2, 16'ha4d2, 16'ha4b2, 16'ha4d2, 16'ha4d2, 16'ha4b2, 16'ha4b1, 16'ha471, 16'h9c30, 16'h9c71, 16'h9c70, 16'h9430, 16'h9450, 16'h9450, 16'h9450, 16'h9c71, 16'h9430, 16'h736d, 16'h9450, 16'ha4d2, 16'ha4d2, 16'ha4d1, 16'ha4b1, 16'h9cb1, 16'h9cb1, 16'h9cb1, 16'h9cb1, 16'h9cb1, 16'h944f, 16'h5aa9, 16'h4a48, 16'h6b4b, 16'h5269, 16'h3165, 16'h5aaa, 16'h4a28, 16'h3985, 16'h3164, 16'h3164, 16'h3144, 16'h2944, 16'h2944, 16'h2944, 16'h2924, 16'h2923, 16'h213, 16'h213, 16'h18c2, 16'h18c2, 16'h5268, 16'h5aa9, 16'h4a27, 16'h2944, 16'h18c2, 16'h4248, 16'h3268, 16'h3227, 16'h427, 16'h18c2, 16'h861, 16'h2944, 16'h5269, 16'h6aeb, 16'h6bb, 16'h5a89, 16'h5aaa, 16'h5aaa, 16'h4a48, 16'h41e7, 16'h41c6, 16'h5289, 16'h6bb, 16'h6b2b, 16'h6bb, 16'h5acb, 16'h5acb, 16'h5aab, 16'h5acb, 16'h6b2b, 16'h6b4c, 16'h6b2b, 16'h6aeb, 16'h62ca, 16'h52aa, 16'h52aa, 16'h52aa, 16'h52aa, 16'h528a, 16'h52aa, 16'h5acb, 16'h62eb, 16'h62ec, 16'h6bb, 16'h6bc, 16'h6b2c, 16'h732c, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h6b2b, 16'h6b2c, 16'h6b2c, 16'h6b2b, 16'h6b2c, 16'h6bb, 16'h63b, 16'h63b, 16'h6bc, 16'h734c, 16'h7b4c, 16'h9c2f, 16'hcdd5, 16'hd5f6, 16'hd5f5, 16'hd5f5, 16'hd5f5, 16'hd5d5, 16'hd5d5, 16'hcdd5, 16'hcdd5, 16'hcdd5, 16'hcdd5, 16'hcdb5, 16'hcdb5, 16'hcdb5, 16'hcdb4, 16'hcdb4, 16'hcd94, 16'hcd94, 16'hcd94, 16'hcd94, 16'hc594, 16'hc594, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc573, 16'hc553, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha44f, 16'ha44f, 16'h7b4b, 16'h3143, 16'h20e2, 16'h20e2, 16'h20c2, 16'h20c2, 16'h1081, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'hb533, 16'hb513, 16'hb4d2, 16'hb513, 16'hb554, 16'hb554, 16'hb513, 16'hb4d2, 16'hb4b2, 16'hb4b2, 16'hacd1, 16'h9c4f, 16'ha490, 16'hacd2, 16'had13, 16'hb533, 16'hacf2, 16'h5aaa, 16'h83ce, 16'h9cb1, 16'ha4d2, 16'ha4d2, 16'h9cb1, 16'h9cb1, 16'h9cb1, 16'h9cb1, 16'h9cb1, 16'ha4d2, 16'ha4f3, 16'h62c9, 16'h3a27, 16'h5aca, 16'h5a89, 16'h4a27, 16'h736c, 16'h5268, 16'h39a5, 16'h3164, 16'h3164, 16'h3164, 16'h2944, 16'h2944, 16'h2924, 16'h2924, 16'h2123, 16'h213, 16'h20e3, 16'h18a2, 16'h213, 16'h5aa9, 16'h5a89, 16'h4a27, 16'h2944, 16'h18c2, 16'h4248, 16'h3248, 16'h3227, 16'h41e7, 16'h18c2, 16'h861, 16'h2944, 16'h5289, 16'h6bb, 16'h6b2b, 16'h5aa9, 16'h5268, 16'h5a89, 16'h4a28, 16'h41e7, 16'h41c6, 16'h5269, 16'h6bb, 16'h6bb, 16'h63b, 16'h5aca, 16'h5acb, 16'h5aab, 16'h5aab, 16'h63b, 16'h6b2b, 16'h6bb, 16'h62eb, 16'h5aca, 16'h52aa, 16'h52aa, 16'h52aa, 16'h52aa, 16'h528a, 16'h52aa, 16'h5acb, 16'h62eb, 16'h62eb, 16'h6bc, 16'h6bc, 16'h6b2c, 16'h6b2c, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h6b4c, 16'h6bb, 16'h6b2b, 16'h6b2c, 16'h6b2b, 16'h6b2b, 16'h6bb, 16'h6bb, 16'h6bb, 16'h6bc, 16'h734c, 16'h734c, 16'h9c4f, 16'hd5f5, 16'hd5f6, 16'hd5f6, 16'hd5f6, 16'hd5f5, 16'hd5f5, 16'hd5d5, 16'hd5d5, 16'hd5d5, 16'hd5d5, 16'hd5d5, 16'hcdd5, 16'hcdd5, 16'hcdd5, 16'hcdb5, 16'hcdb5, 16'hcdb5, 16'hcdb4, 16'hcd94, 16'hcd94, 16'hcd94, 16'hcd94, 16'hc594, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc573, 16'hc573, 16'hc573, 16'hc553, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha44f, 16'h7b4b, 16'h3144, 16'h20e2, 16'h20e2, 16'h20e2, 16'h20c2, 16'h1061, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'hb513, 16'hb4f3, 16'hbcf3, 16'hb513, 16'hb533, 16'hb533, 16'hb533, 16'hb513, 16'hb533, 16'hb4f2, 16'hb4d2, 16'hac50, 16'hac50, 16'hb492, 16'had13, 16'hb533, 16'ha4d2, 16'h5aa9, 16'h83ce, 16'h9cb1, 16'ha4d2, 16'ha4d1, 16'ha4b1, 16'h9cb1, 16'h9cb1, 16'h9cb1, 16'ha4b1, 16'hb534, 16'hc5d6, 16'h6ba, 16'h31c6, 16'h4a48, 16'h41e7, 16'h5289, 16'h944f, 16'h5aa9, 16'h39a6, 16'h3185, 16'h3164, 16'h3164, 16'h2944, 16'h2944, 16'h2944, 16'h2924, 16'h213, 16'h213, 16'h18c2, 16'h1081, 16'h39a6, 16'h62ca, 16'h5a89, 16'h4a7, 16'h2944, 16'h20e3, 16'h4a68, 16'h3228, 16'h3227, 16'h39e7, 16'h10a2, 16'h861, 16'h2944, 16'h5a89, 16'h6b2b, 16'h6b2b, 16'h62ea, 16'h5248, 16'h4a28, 16'h41e7, 16'h41e7, 16'h39c6, 16'h5268, 16'h62ea, 16'h62ea, 16'h63b, 16'h5aca, 16'h5aca, 16'h5aaa, 16'h5aaa, 16'h62eb, 16'h6aeb, 16'h6bb, 16'h62eb, 16'h5aca, 16'h528a, 16'h52aa, 16'h52aa, 16'h528a, 16'h528a, 16'h52aa, 16'h5acb, 16'h62cb, 16'h62eb, 16'h6bc, 16'h6bc, 16'h6bb, 16'h6b2b, 16'h732b, 16'h734c, 16'h734c, 16'h734c, 16'h734c, 16'h6b4c, 16'h6b2b, 16'h6b2b, 16'h6b2b, 16'h6b2b, 16'h6b2c, 16'h6b2b, 16'h6bb, 16'h6aeb, 16'h6bb, 16'h734c, 16'h736c, 16'h9c50, 16'hd5f6, 16'hd616, 16'hd616, 16'hd616, 16'hd5f6, 16'hd5f6, 16'hd5f5, 16'hd5f5, 16'hd5f5, 16'hd5f5, 16'hd5d5, 16'hd5d5, 16'hd5d5, 16'hcdd5, 16'hcdd5, 16'hcdd5, 16'hcdb5, 16'hcdb5, 16'hcdb4, 16'hcdb4, 16'hcdb4, 16'hcd94, 16'hcd94, 16'hc594, 16'hc594, 16'hc594, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc573, 16'hc573, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha44f, 16'h7b4b, 16'h3144, 16'h20e2, 16'h20e2, 16'h20e2, 16'h20e2, 16'h1081, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'hb4f3, 16'hb513, 16'hb513, 16'hb513, 16'hb513, 16'hb513, 16'hb513, 16'hb513, 16'hb513, 16'hb4d2, 16'hb4d2, 16'hb4b1, 16'hb471, 16'hac91, 16'hacf2, 16'hb533, 16'ha4d1, 16'h5aa9, 16'h83cd, 16'h9cb1, 16'ha4d2, 16'ha4b2, 16'ha4b2, 16'h9cb1, 16'h9cb1, 16'h9cb1, 16'ha4f2, 16'hbd95, 16'hbdb5, 16'h62a9, 16'h2965, 16'h4a28, 16'h41c6, 16'h6b2b, 16'h9c90, 16'h736c, 16'h41c6, 16'h3185, 16'h3165, 16'h3164, 16'h2944, 16'h2944, 16'h2924, 16'h213, 16'h18e3, 16'h18c2, 16'h10a2, 16'h1081, 16'h41c6, 16'h62a9, 16'h5268, 16'h4a7, 16'h2944, 16'h213, 16'h4268, 16'h2a27, 16'h29e6, 16'h2985, 16'h1081, 16'h841, 16'h2124, 16'h5269, 16'h6bb, 16'h6b2b, 16'h62ca, 16'h4a48, 16'h3985, 16'h3185, 16'h41e7, 16'h41c6, 16'h5268, 16'h62eb, 16'h62ea, 16'h63b, 16'h5aca, 16'h5aaa, 16'h52aa, 16'h5aaa, 16'h62ca, 16'h62ea, 16'h62ea, 16'h62ea, 16'h5aca, 16'h5289, 16'h528a, 16'h52aa, 16'h528a, 16'h528a, 16'h52aa, 16'h5acb, 16'h62cb, 16'h62eb, 16'h6bc, 16'h6bc, 16'h6bb, 16'h6b2b, 16'h732c, 16'h734c, 16'h732c, 16'h6b2c, 16'h734c, 16'h734c, 16'h6b2b, 16'h6b2b, 16'h6bb, 16'h6bc, 16'h6b2c, 16'h6bb, 16'h6bb, 16'h62eb, 16'h6bb, 16'h734c, 16'h736c, 16'h9c50, 16'hd616, 16'hd636, 16'hd616, 16'hd616, 16'hd616, 16'hd616, 16'hd616, 16'hd5f6, 16'hd5f6, 16'hd5f6, 16'hd5f6, 16'hd5d5, 16'hd5d5, 16'hd5d5, 16'hd5d5, 16'hd5d5, 16'hd5d5, 16'hcdd5, 16'hcdb5, 16'hcdb5, 16'hcdb5, 16'hcdb4, 16'hcd94, 16'hcd94, 16'hcd94, 16'hc594, 16'hc594, 16'hc594, 16'hc574, 16'hc574, 16'hc574, 16'hc573, 16'hc573, 16'hc553, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'h836b, 16'h3143, 16'h20e2, 16'h20e2, 16'h20e2, 16'h20e2, 16'h1081, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'hbcf3, 16'hbcf3, 16'hbcf3, 16'hb513, 16'hb513, 16'hb513, 16'hb4f3, 16'hb4d2, 16'hb4d2, 16'hb4d2, 16'hb4f2, 16'hacd2, 16'hb491, 16'hac91, 16'hacf2, 16'hb533, 16'ha4b1, 16'h5a89, 16'h83ad, 16'h9cb1, 16'ha4d2, 16'h9470, 16'h9450, 16'h9cb1, 16'ha4b1, 16'ha4b1, 16'ha4d2, 16'had13, 16'ha4d2, 16'h5a89, 16'h31c6, 16'h39e7, 16'h39a6, 16'h6bb, 16'h736c, 16'h6b2b, 16'h427, 16'h3165, 16'h3164, 16'h2944, 16'h2944, 16'h2944, 16'h213, 16'h18c3, 16'h10a2, 16'h1082, 16'h861, 16'h841, 16'h18c2, 16'h4a27, 16'h5248, 16'h427, 16'h3144, 16'h20e3, 16'h2985, 16'h2185, 16'h113, 16'h861, 16'h840, 16'h840, 16'h18a2, 16'h3185, 16'h41c6, 16'h41e6, 16'h39a6, 16'h3185, 16'h3185, 16'h39c6, 16'h39c6, 16'h39a6, 16'h5269, 16'h63b, 16'h6b2b, 16'h6b2b, 16'h62eb, 16'h5acb, 16'h5aaa, 16'h5aaa, 16'h62ca, 16'h62ca, 16'h62ca, 16'h62ca, 16'h5aca, 16'h528a, 16'h528a, 16'h528a, 16'h528a, 16'h528a, 16'h5aaa, 16'h5acb, 16'h62eb, 16'h63b, 16'h6bb, 16'h6bb, 16'h6bb, 16'h6b2b, 16'h6b2c, 16'h732c, 16'h6b2b, 16'h6b2b, 16'h6b2c, 16'h6b2c, 16'h6b2b, 16'h6b2b, 16'h6bb, 16'h6bb, 16'h6b2b, 16'h6bb, 16'h6bb, 16'h62eb, 16'h6bb, 16'h734c, 16'h734c, 16'h9c50, 16'hd636, 16'hde36, 16'hde36, 16'hd616, 16'hde16, 16'hd616, 16'hd616, 16'hd616, 16'hd616, 16'hd5f6, 16'hd5f6, 16'hd5f6, 16'hd5f6, 16'hd5f5, 16'hd5d5, 16'hd5d5, 16'hd5d5, 16'hd5d5, 16'hcdd5, 16'hcdd5, 16'hcdb5, 16'hcdb5, 16'hcdb4, 16'hcdb4, 16'hcdb4, 16'hcd94, 16'hcd94, 16'hc594, 16'hc594, 16'hc594, 16'hc574, 16'hc574, 16'hc573, 16'hc573, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4d2, 16'hacd1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'h836b, 16'h3143, 16'h20e2, 16'h20e2, 16'h20e2, 16'h20c2, 16'h1081, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'hbcd3, 16'hbcf3, 16'hbd13, 16'hb513, 16'hb533, 16'had13, 16'hb513, 16'hb4f2, 16'hb4b2, 16'hb492, 16'had13, 16'hacf2, 16'hacf2, 16'hacf2, 16'had12, 16'hb533, 16'h9cb1, 16'h5a89, 16'h83cd, 16'h9cb1, 16'h9cb1, 16'h7bad, 16'h5a89, 16'h7bae, 16'ha4b1, 16'ha4b1, 16'ha4b1, 16'h9c70, 16'h944f, 16'h62ea, 16'h29e6, 16'h31c6, 16'h2965, 16'h2965, 16'h2965, 16'h2965, 16'h2965, 16'h3185, 16'h39c6, 16'h31a5, 16'h213, 16'h2123, 16'h10a2, 16'h1061, 16'h1082, 16'h861, 16'h861, 16'h841, 16'h10a2, 16'h41e6, 16'h4a27, 16'h41c6, 16'h2944, 16'h1081, 16'h8a1, 16'h8a2, 16'h881, 16'h840, 16'h840, 16'h840, 16'h841, 16'h20e3, 16'h2944, 16'h3165, 16'h2924, 16'h2124, 16'h20e3, 16'h213, 16'h2944, 16'h3986, 16'h5268, 16'h6bb, 16'h6b2b, 16'h6b2c, 16'h734c, 16'h6b2b, 16'h62eb, 16'h62ca, 16'h62ca, 16'h62ca, 16'h62ea, 16'h62ca, 16'h5aca, 16'h528a, 16'h528a, 16'h528a, 16'h528a, 16'h528a, 16'h5aaa, 16'h62cb, 16'h62eb, 16'h6bb, 16'h6bc, 16'h6b2c, 16'h6b2c, 16'h6b2c, 16'h6b2b, 16'h6b2c, 16'h6bc, 16'h6b2c, 16'h6b2c, 16'h6b2c, 16'h6bb, 16'h6bb, 16'h6bb, 16'h6b2b, 16'h6b2b, 16'h6b2b, 16'h6bb, 16'h62eb, 16'h6bb, 16'h734c, 16'h734c, 16'h9c50, 16'hde37, 16'hde57, 16'hde57, 16'hde36, 16'hde36, 16'hde36, 16'hd636, 16'hd616, 16'hd616, 16'hd616, 16'hd616, 16'hd5f6, 16'hd5f6, 16'hd5f6, 16'hd5f6, 16'hd5f5, 16'hd5d5, 16'hd5d5, 16'hd5d5, 16'hd5d5, 16'hcdd5, 16'hcdd5, 16'hcdb5, 16'hcdb5, 16'hcdb5, 16'hcdb4, 16'hcdb4, 16'hcd94, 16'hcd94, 16'hcd94, 16'hc594, 16'hc594, 16'hc574, 16'hc573, 16'hc573, 16'hc553, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4d2, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'h836b, 16'h3143, 16'h20e2, 16'h20e2, 16'h20e2, 16'h20c2, 16'h1081, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'hbcd2, 16'hb4f3, 16'hb4f3, 16'hb4d2, 16'hb513, 16'had13, 16'had13, 16'hb513, 16'hb4f3, 16'hb4f3, 16'had13, 16'hacd2, 16'hacf2, 16'hacf2, 16'had12, 16'hb533, 16'h9c90, 16'h5a89, 16'h83ad, 16'h9cb1, 16'h8cf, 16'h4a28, 16'h18c3, 16'h3165, 16'h736c, 16'ha4b1, 16'ha4b1, 16'h9c91, 16'h942f, 16'h6bb, 16'h327, 16'h4aaa, 16'h6b4c, 16'h52ca, 16'h4a69, 16'h4a69, 16'h4a69, 16'h4268, 16'h4268, 16'h3a27, 16'h2165, 16'h29a6, 16'h2965, 16'h20e3, 16'h2124, 16'h214, 16'h214, 16'h2124, 16'h2124, 16'h2965, 16'h2964, 16'h2924, 16'h18c2, 16'h10a2, 16'h1944, 16'h1944, 16'h1924, 16'h18e2, 16'h18c2, 16'h1081, 16'h18a2, 16'h427, 16'h62ca, 16'h62ea, 16'h5269, 16'h4a68, 16'h39a6, 16'h2124, 16'h20e3, 16'h2924, 16'h4a48, 16'h6bb, 16'h6b2b, 16'h6b2c, 16'h734c, 16'h732c, 16'h6b2b, 16'h6bb, 16'h6b2b, 16'h6bb, 16'h6aea, 16'h62ea, 16'h62ca, 16'h5289, 16'h5289, 16'h5289, 16'h528a, 16'h528a, 16'h5aaa, 16'h5acb, 16'h62eb, 16'h62eb, 16'h6b2c, 16'h6b2c, 16'h6b2c, 16'h6b2b, 16'h6b2b, 16'h6b2c, 16'h6b2b, 16'h6b2b, 16'h6b2b, 16'h6b2b, 16'h6bb, 16'h6bb, 16'h6bb, 16'h6b2b, 16'h6bb, 16'h6bb, 16'h6bb, 16'h62eb, 16'h6bb, 16'h732c, 16'h734c, 16'h9c70, 16'hde57, 16'hde77, 16'hde77, 16'hde57, 16'hde57, 16'hde37, 16'hde36, 16'hde36, 16'hde36, 16'hde36, 16'hd616, 16'hd616, 16'hd616, 16'hd5f6, 16'hd5f6, 16'hd5f6, 16'hd5f6, 16'hd5f5, 16'hd5f5, 16'hd5d5, 16'hd5d5, 16'hcdd5, 16'hcdd5, 16'hcdd5, 16'hcdb5, 16'hcdb5, 16'hcdb4, 16'hcdb4, 16'hcd94, 16'hcd94, 16'hcd94, 16'hc594, 16'hc574, 16'hc574, 16'hc574, 16'hc573, 16'hc573, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'h836c, 16'h3144, 16'h28e2, 16'h20e2, 16'h20c2, 16'h20c2, 16'h1081, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'hb4d3, 16'hb4f2, 16'hb4b2, 16'hb492, 16'hacf2, 16'had12, 16'had33, 16'hb533, 16'hb533, 16'had33, 16'had13, 16'hacf2, 16'hacf2, 16'hacf2, 16'had12, 16'hb512, 16'h9c70, 16'h5a69, 16'h7b8d, 16'h83ce, 16'h41e7, 16'h10a2, 16'h1081, 16'h1081, 16'h214, 16'h62ea, 16'h9c70, 16'ha4b2, 16'ha4b1, 16'h83ce, 16'h4a89, 16'h4a68, 16'h4aa9, 16'h4aa9, 16'h3a27, 16'h31e6, 16'h31c6, 16'h31e6, 16'h31c6, 16'h29a6, 16'h29a5, 16'h29c5, 16'h39e6, 16'h3185, 16'h213, 16'h18a2, 16'h1082, 16'h1082, 16'h1082, 16'h1082, 16'h1061, 16'h1061, 16'h861, 16'h841, 16'h861, 16'h861, 16'h861, 16'h861, 16'h861, 16'h840, 16'h861, 16'h18c2, 16'h20e3, 16'h213, 16'h18c2, 16'h18e3, 16'h18c2, 16'h10a2, 16'h1081, 16'h1081, 16'h41c6, 16'h63b, 16'h6bb, 16'h732c, 16'h734c, 16'h6b2b, 16'h6bb, 16'h6b2b, 16'h734c, 16'h736c, 16'h6bb, 16'h6aeb, 16'h62ea, 16'h5aaa, 16'h5aaa, 16'h5289, 16'h528a, 16'h528a, 16'h52aa, 16'h5acb, 16'h62cb, 16'h62eb, 16'h6bc, 16'h6b2c, 16'h6b2c, 16'h6b2b, 16'h6b2b, 16'h6bb, 16'h6b2b, 16'h6b2b, 16'h6b2b, 16'h6b2b, 16'h6bb, 16'h6bb, 16'h6bb, 16'h6bb, 16'h6bb, 16'h6bb, 16'h6aeb, 16'h62eb, 16'h6aeb, 16'h732b, 16'h734c, 16'h9c70, 16'hde77, 16'he678, 16'he678, 16'hde77, 16'hde57, 16'hde57, 16'hde57, 16'hde37, 16'hde36, 16'hde36, 16'hde36, 16'hd636, 16'hd616, 16'hd616, 16'hd616, 16'hd616, 16'hd5f6, 16'hd5f6, 16'hd5f6, 16'hd5f6, 16'hd5f5, 16'hd5d5, 16'hd5d5, 16'hcdd5, 16'hcdd5, 16'hcdb5, 16'hcdb5, 16'hcdb4, 16'hcdb4, 16'hcd94, 16'hcd94, 16'hc594, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc553, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'h836c, 16'h3144, 16'h20e2, 16'h20e2, 16'h20c2, 16'h20e2, 16'h1081, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'hb4b2, 16'hb4f2, 16'hb4b2, 16'hb471, 16'hacd2, 16'had12, 16'had12, 16'had13, 16'had13, 16'hb533, 16'hb513, 16'hacd2, 16'hacf2, 16'hacf2, 16'hacf2, 16'had12, 16'h83ad, 16'h3145, 16'h5269, 16'h5aca, 16'h39c6, 16'h18a2, 16'h1081, 16'h1061, 16'h1082, 16'h3986, 16'h7b6d, 16'ha4b1, 16'ha4d2, 16'ha4b1, 16'h83ac, 16'h6ac9, 16'h6ae9, 16'h6ba, 16'h5268, 16'h3165, 16'h3165, 16'h3164, 16'h3164, 16'h2944, 16'h2944, 16'h2943, 16'h2924, 16'h293, 16'h20c3, 16'h18a2, 16'h18a2, 16'h1082, 16'h1082, 16'h1081, 16'h1061, 16'h861, 16'h840, 16'h840, 16'h820, 16'h840, 16'h861, 16'h841, 16'h840, 16'h840, 16'h18c2, 16'h39a6, 16'h4a28, 16'h4a28, 16'h41c6, 16'h3165, 16'h2944, 16'h2965, 16'h39a6, 16'h39c6, 16'h5aa9, 16'h6b2b, 16'h6b2b, 16'h6bb, 16'h6bb, 16'h6aea, 16'h6aea, 16'h6b2b, 16'h6bb, 16'h736c, 16'h6b2b, 16'h6b2b, 16'h6bb, 16'h6bb, 16'h6bb, 16'h734b, 16'h83ad, 16'h62ea, 16'h5289, 16'h5aca, 16'h62eb, 16'h62eb, 16'h6bb, 16'h6b2c, 16'h6b2b, 16'h6b2b, 16'h6b2b, 16'h6bb, 16'h6b2b, 16'h6b2b, 16'h6b2b, 16'h6bb, 16'h6bb, 16'h6ba, 16'h6bb, 16'h6bb, 16'h6bb, 16'h6bb, 16'h62eb, 16'h62ca, 16'h62ea, 16'h732b, 16'h732b, 16'h9c50, 16'he678, 16'he698, 16'he698, 16'he678, 16'he677, 16'hde77, 16'hde57, 16'hde57, 16'hde37, 16'hde37, 16'hde36, 16'hd636, 16'hd636, 16'hd616, 16'hd616, 16'hd616, 16'hd616, 16'hd616, 16'hd5f6, 16'hd5f6, 16'hd5f6, 16'hd5d5, 16'hd5d5, 16'hd5d5, 16'hd5d5, 16'hcdd5, 16'hcdb5, 16'hcdb5, 16'hcdb5, 16'hcdb4, 16'hcd94, 16'hcd94, 16'hc594, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc573, 16'hc573, 16'hc573, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd12, 16'hbd12, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb1, 16'hacb1, 16'ha4b0, 16'hacb0, 16'hac90, 16'hac90, 16'ha490, 16'ha470, 16'h836b, 16'h3143, 16'h212, 16'h20e2, 16'h20e2, 16'h20e2, 16'h1081, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'hb4f2, 16'hb512, 16'hb4f2, 16'hacb1, 16'hacf2, 16'had12, 16'had12, 16'had12, 16'hacf2, 16'hacd2, 16'hacd2, 16'hacd2, 16'hacf2, 16'hacf2, 16'hacf2, 16'had12, 16'h7b6c, 16'h2944, 16'h5a89, 16'h7b6d, 16'h83ce, 16'h62ca, 16'h39a5, 16'h20e3, 16'h5248, 16'h8c2f, 16'ha4d1, 16'had13, 16'hacf2, 16'ha4d1, 16'h8bed, 16'h73a, 16'h6ae9, 16'h739, 16'h5a88, 16'h1882, 16'h1062, 16'h1882, 16'h1041, 16'h1041, 16'h841, 16'h841, 16'h841, 16'h1041, 16'h1041, 16'h1061, 16'h1061, 16'h1061, 16'h1061, 16'h1061, 16'h1061, 16'h1061, 16'h861, 16'h1061, 16'h1061, 16'h1081, 16'h18e2, 16'h18a2, 16'h1061, 16'h1061, 16'h213, 16'h4a7, 16'h5a68, 16'h5a88, 16'h5248, 16'h4a7, 16'h41e6, 16'h4a7, 16'h5269, 16'h5269, 16'h62ea, 16'h736c, 16'h736c, 16'h734c, 16'h732b, 16'h734b, 16'h7b4b, 16'h7b6b, 16'h7b6b, 16'h7b6c, 16'h732b, 16'h836b, 16'h838c, 16'h7b4b, 16'h6ae9, 16'h6ac8, 16'h6ac9, 16'h5226, 16'h5247, 16'h62aa, 16'h62ca, 16'h62ea, 16'h6aea, 16'h6aea, 16'h6aea, 16'h6aea, 16'h6aea, 16'h62ea, 16'h6aea, 16'h6aea, 16'h62ea, 16'h62ea, 16'h62ea, 16'h62ea, 16'h62ea, 16'h62ea, 16'h6aea, 16'h6aea, 16'h6aea, 16'h6aea, 16'h6aea, 16'h6aea, 16'h6ba, 16'h9c4f, 16'hee98, 16'hee98, 16'he698, 16'he698, 16'he678, 16'he677, 16'hde57, 16'hde57, 16'hde57, 16'hde57, 16'hde37, 16'hde37, 16'hde36, 16'hde36, 16'hd636, 16'hd636, 16'hd616, 16'hd616, 16'hd616, 16'hd616, 16'hd5f6, 16'hd5f5, 16'hd5f5, 16'hd5d5, 16'hd5d5, 16'hcdd5, 16'hcdd5, 16'hcdb5, 16'hcdb5, 16'hcdb4, 16'hcdb4, 16'hcd94, 16'hcd94, 16'hc594, 16'hc594, 16'hc574, 16'hc574, 16'hc574, 16'hc573, 16'hc573, 16'hc553, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f2, 16'hb4d1, 16'hb4d2, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hac90, 16'ha490, 16'ha490, 16'h836c, 16'h3143, 16'h20e2, 16'h20e2, 16'h20e2, 16'h20c2, 16'h1081, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'hb513, 16'hb533, 16'hb533, 16'had12, 16'had12, 16'had32, 16'had12, 16'had12, 16'hacd2, 16'hac91, 16'hacb1, 16'hacd2, 16'ha4d2, 16'ha4d2, 16'hacf2, 16'had13, 16'h944f, 16'h5268, 16'h6b2b, 16'h7b8d, 16'h734d, 16'h732b, 16'h5a89, 16'h4a7, 16'h62ea, 16'h734c, 16'h83ae, 16'hbd74, 16'hb533, 16'hacd1, 16'h8bed, 16'h73a, 16'h73a, 16'h732a, 16'h6288, 16'h1882, 16'h3145, 16'h6b2b, 16'h41c6, 16'h20e3, 16'h18c2, 16'h18c3, 16'h214, 16'h3145, 16'h3185, 16'h3985, 16'h3985, 16'h3985, 16'h3165, 16'h3144, 16'h2924, 16'h213, 16'h213, 16'h2124, 16'h214, 16'h193, 16'h213, 16'h18e2, 16'h18a2, 16'h10a2, 16'h20e2, 16'h3164, 16'h41a5, 16'h41c6, 16'h39a5, 16'h3984, 16'h3984, 16'h41c6, 16'h4a27, 16'h4a48, 16'h62ea, 16'h736c, 16'h736c, 16'h736c, 16'h8bcd, 16'h9c6f, 16'h93ed, 16'h8bcd, 16'h7b4b, 16'h6aea, 16'h6aea, 16'h6ae9, 16'h5a47, 16'h49e5, 16'h41c5, 16'h3984, 16'h3163, 16'h3123, 16'h41a5, 16'h5268, 16'h62a9, 16'h62c9, 16'h62c9, 16'h62c9, 16'h62c9, 16'h62c9, 16'h62c9, 16'h62c9, 16'h62c9, 16'h62c9, 16'h62c9, 16'h62c9, 16'h62c9, 16'h62ca, 16'h62ca, 16'h62ca, 16'h6aca, 16'h6aca, 16'h6aca, 16'h6aea, 16'h6aea, 16'h6aea, 16'h6aea, 16'h9c4f, 16'hee98, 16'heeb9, 16'heeb8, 16'he698, 16'he698, 16'he678, 16'he677, 16'hde77, 16'hde57, 16'hde57, 16'hde57, 16'hde57, 16'hde37, 16'hde36, 16'hde36, 16'hde36, 16'hd636, 16'hd616, 16'hd616, 16'hd616, 16'hd5f6, 16'hd5f6, 16'hd5f5, 16'hd5f5, 16'hd5d5, 16'hd5d5, 16'hcdd5, 16'hcdb5, 16'hcdb5, 16'hcdb5, 16'hcdb4, 16'hcdb4, 16'hcd94, 16'hc594, 16'hc594, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc573, 16'hc553, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'ha490, 16'ha490, 16'h836c, 16'h3144, 16'h20e3, 16'h20e2, 16'h20e2, 16'h20c2, 16'h1081, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'hb533, 16'hb553, 16'hb533, 16'had33, 16'hb533, 16'had32, 16'had12, 16'had12, 16'hacd2, 16'hacb1, 16'hacb1, 16'hacb2, 16'hacf2, 16'hacf2, 16'hacf2, 16'had12, 16'h9450, 16'h5a89, 16'h83ce, 16'ha4d2, 16'hacf2, 16'ha4d2, 16'h9cb1, 16'h9450, 16'h7b8c, 16'h4a7, 16'h62ca, 16'hb533, 16'hacf2, 16'h9c50, 16'h8bad, 16'h73a, 16'h73a, 16'h732a, 16'h62a8, 16'h1882, 16'h4165, 16'ha4b0, 16'h942e, 16'h4a47, 16'h2923, 16'h2124, 16'h3165, 16'h39a6, 16'h41c6, 16'h41c6, 16'h41c6, 16'h41a6, 16'h39a5, 16'h3185, 16'h2944, 16'h2944, 16'h2944, 16'h2944, 16'h2944, 16'h2944, 16'h2923, 16'h2923, 16'h213, 16'h293, 16'h2944, 16'h3984, 16'h41c5, 16'h41c6, 16'h3144, 16'h28e2, 16'h28e2, 16'h28e2, 16'h313, 16'h3943, 16'h5a68, 16'h6b4c, 16'h734c, 16'h7b6d, 16'h9c4f, 16'h94d, 16'h739, 16'h9c2e, 16'h9c4f, 16'h9c2e, 16'h93ed, 16'h6ac9, 16'h526, 16'h5a47, 16'h4a7, 16'h3144, 16'h20c2, 16'h20e3, 16'h3985, 16'h5247, 16'h5a89, 16'h62a9, 16'h62a9, 16'h62a9, 16'h62a9, 16'h62a9, 16'h62a9, 16'h62c9, 16'h62c9, 16'h62a9, 16'h62a9, 16'h62a9, 16'h62c9, 16'h62a9, 16'h62a9, 16'h62c9, 16'h62c9, 16'h62c9, 16'h62c9, 16'h62c9, 16'h62c9, 16'h6ac9, 16'h6aca, 16'h9c2f, 16'heeb8, 16'heeb9, 16'heeb9, 16'heeb8, 16'he698, 16'he678, 16'he678, 16'hde77, 16'hde77, 16'hde57, 16'hde57, 16'hde57, 16'hde37, 16'hde36, 16'hde36, 16'hde36, 16'hde36, 16'hd636, 16'hd616, 16'hd616, 16'hd616, 16'hd5f5, 16'hd5f5, 16'hd5f5, 16'hd5f5, 16'hd5d5, 16'hcdd5, 16'hcdd5, 16'hcdb5, 16'hcdb5, 16'hcdb5, 16'hcdb4, 16'hcd94, 16'hcd94, 16'hc594, 16'hc594, 16'hc574, 16'hc574, 16'hc574, 16'hc573, 16'hc573, 16'hc553, 16'hc553, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4d1, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'ha4b1, 16'hacb1, 16'ha490, 16'h838c, 16'h3143, 16'h20e2, 16'h20e2, 16'h20e2, 16'h20c2, 16'h1081, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'had12, 16'had33, 16'hb533, 16'had33, 16'hb533, 16'hb533, 16'had12, 16'had13, 16'hacf2, 16'hacd2, 16'hacd2, 16'hacb2, 16'hacf2, 16'had12, 16'hacf2, 16'had12, 16'h9c6f, 16'h5a89, 16'h8bee, 16'ha4d2, 16'hacf2, 16'hacf2, 16'hacf2, 16'hacf2, 16'hacf2, 16'h734c, 16'h732c, 16'hb533, 16'hbd95, 16'ha4d2, 16'h83ad, 16'h73a, 16'h73a, 16'h7b2b, 16'h734a, 16'h5227, 16'h6269, 16'h8bad, 16'h94e, 16'h736b, 16'h39a4, 16'h39a5, 16'h41e6, 16'h4a6, 16'h4a6, 16'h4a6, 16'h49e6, 16'h49e6, 16'h41c6, 16'h41c6, 16'h41c5, 16'h41a5, 16'h39a5, 16'h39a5, 16'h39c5, 16'h41c5, 16'h41c6, 16'h41c6, 16'h41c6, 16'h41c6, 16'h49e6, 16'h5a47, 16'h5247, 16'h4a6, 16'h3144, 16'h3124, 16'h3144, 16'h3164, 16'h3964, 16'h4185, 16'h5a89, 16'h734c, 16'h7b8d, 16'h83ad, 16'hacb0, 16'h94d, 16'h6aa8, 16'h8bcd, 16'h8bcd, 16'h93ed, 16'h94d, 16'h94d, 16'h93ed, 16'h83ac, 16'h6aea, 16'h5247, 16'h4a6, 16'h4a7, 16'h5247, 16'h5a88, 16'h62a9, 16'h62a9, 16'h62a9, 16'h5a88, 16'h5aa8, 16'h62a8, 16'h62a8, 16'h62a8, 16'h62a8, 16'h62a8, 16'h6288, 16'h62a8, 16'h62a8, 16'h62a8, 16'h62a8, 16'h62a8, 16'h62a9, 16'h62a9, 16'h6288, 16'h6288, 16'h6288, 16'h62a8, 16'h62a9, 16'h94e, 16'heeb8, 16'heeb9, 16'heeb9, 16'heeb9, 16'hee98, 16'he698, 16'he698, 16'he678, 16'he678, 16'hde77, 16'hde57, 16'hde57, 16'hde57, 16'hde37, 16'hde37, 16'hde36, 16'hde36, 16'hde36, 16'hd616, 16'hd616, 16'hd616, 16'hd5f6, 16'hd5f5, 16'hd5f6, 16'hd5f5, 16'hd5d5, 16'hcdd5, 16'hcdd5, 16'hcdb5, 16'hcdb5, 16'hcdb5, 16'hcdb4, 16'hcd94, 16'hcd94, 16'hc594, 16'hc594, 16'hc594, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc573, 16'hc553, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd32, 16'hbd33, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'ha490, 16'h838c, 16'h3164, 16'h20e2, 16'h20e2, 16'h20e2, 16'h20e2, 16'h1081, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'hb4f2, 16'hb513, 16'hb513, 16'hb533, 16'hb533, 16'hb533, 16'hb532, 16'hb533, 16'hb533, 16'hb4d2, 16'hacf2, 16'hacf2, 16'had12, 16'had12, 16'had12, 16'had32, 16'h9c6f, 16'h5a89, 16'h8bee, 16'ha4d2, 16'had12, 16'had12, 16'hacf2, 16'h8bef, 16'h8bef, 16'h7b6c, 16'h6aa9, 16'ha490, 16'hbd54, 16'h7b6e, 16'h628a, 16'h73a, 16'h6ac9, 16'h7b2b, 16'h7b4b, 16'h7b2b, 16'h732b, 16'h7b4b, 16'h838c, 16'h736b, 16'h293, 16'h18a2, 16'h18a2, 16'h1882, 16'h1882, 16'h1082, 16'h1061, 16'h1061, 16'h1061, 16'h1061, 16'h1061, 16'h1041, 16'h20c3, 16'h41c7, 16'h4a7, 16'h5248, 16'h5a69, 16'h5a89, 16'h62a9, 16'h62a9, 16'h6aca, 16'h6aea, 16'h6ae9, 16'h6aea, 16'h6aea, 16'h6aeb, 16'h6bb, 16'h6ba, 16'h73a, 16'h73a, 16'h73b, 16'h732b, 16'h7b4c, 16'h838c, 16'h8bcd, 16'h7b4b, 16'h6268, 16'h6288, 16'h41c6, 16'h4a6, 16'h5a68, 16'h526, 16'h5a88, 16'h6ae9, 16'h6ac9, 16'h5268, 16'h41e6, 16'h4a6, 16'h4a6, 16'h4a6, 16'h4a6, 16'h4a26, 16'h4a26, 16'h4a6, 16'h4a6, 16'h4a6, 16'h4a6, 16'h4a6, 16'h4a6, 16'h4a6, 16'h4a6, 16'h4a6, 16'h4a6, 16'h4a6, 16'h4a6, 16'h4a6, 16'h49e6, 16'h49e6, 16'h49e6, 16'h49e5, 16'h49e5, 16'h4a6, 16'h4a6, 16'h8bad, 16'hee98, 16'heeb8, 16'heeb9, 16'heeb9, 16'heeb8, 16'he698, 16'he698, 16'he698, 16'he698, 16'he678, 16'hde77, 16'hde57, 16'hde57, 16'hde57, 16'hde57, 16'hde57, 16'hde57, 16'hde37, 16'hde36, 16'hde16, 16'hd616, 16'hd5f6, 16'hd5f6, 16'hd5f5, 16'hd5f5, 16'hd5f5, 16'hd5d5, 16'hd5d5, 16'hcdb5, 16'hcdb5, 16'hcdb5, 16'hcdb4, 16'hcd94, 16'hcd94, 16'hcd94, 16'hcd94, 16'hc594, 16'hc594, 16'hc594, 16'hc574, 16'hc574, 16'hc573, 16'hc573, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4d1, 16'hb4f1, 16'hb4d1, 16'hacd1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'ha490, 16'h838c, 16'h3164, 16'h212, 16'h20e2, 16'h20e2, 16'h20e2, 16'h1081, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'hacd2, 16'hacf2, 16'hb4f2, 16'hb4f3, 16'hb513, 16'hb533, 16'hb533, 16'hb533, 16'hb533, 16'hb4d2, 16'hb512, 16'hb512, 16'had12, 16'hb512, 16'had12, 16'hb533, 16'h9c6f, 16'h5a89, 16'h8bee, 16'hacf2, 16'had12, 16'had12, 16'had12, 16'h9430, 16'h94f, 16'h8bee, 16'h73b, 16'h7b8c, 16'h7b8d, 16'h4a9, 16'h3966, 16'h7b6c, 16'h7b8d, 16'h83ae, 16'h83ad, 16'h7b4b, 16'h7b4b, 16'h7b4b, 16'h838c, 16'h7b6b, 16'h20e2, 16'h841, 16'h841, 16'h841, 16'h841, 16'h841, 16'h841, 16'h841, 16'h840, 16'h840, 16'h841, 16'h1041, 16'h5248, 16'h83ee, 16'h5a68, 16'h5a68, 16'h5a89, 16'h5aaa, 16'h5a89, 16'h62a9, 16'h6aea, 16'h6289, 16'h5a48, 16'h5248, 16'h5248, 16'h5248, 16'h5248, 16'h5248, 16'h5227, 16'h4a7, 16'h527, 16'h4a7, 16'h4a7, 16'h4a7, 16'h527, 16'h4a6, 16'h41c5, 16'h3985, 16'h213, 16'h18c2, 16'h2923, 16'h18c2, 16'h18a1, 16'h1061, 16'h841, 16'h841, 16'h1081, 16'h3143, 16'h3123, 16'h3163, 16'h3984, 16'h3984, 16'h3143, 16'h3964, 16'h3984, 16'h41a5, 16'h41a5, 16'h41a5, 16'h41c5, 16'h41c5, 16'h41c5, 16'h41c5, 16'h41c5, 16'h41c5, 16'h41c5, 16'h41c5, 16'h41c5, 16'h41c5, 16'h41c5, 16'h41c5, 16'h41e5, 16'h41e5, 16'h49e6, 16'h83ad, 16'hee98, 16'heeb9, 16'heeb9, 16'heeb9, 16'hee98, 16'he698, 16'he698, 16'he698, 16'he678, 16'he678, 16'hde77, 16'hde57, 16'hde57, 16'hde57, 16'hde57, 16'hde57, 16'hde57, 16'hde37, 16'hde36, 16'hde16, 16'hd616, 16'hd5f6, 16'hd5f6, 16'hd5f6, 16'hd5f6, 16'hd5f5, 16'hd5d5, 16'hd5d5, 16'hcdb5, 16'hcdb5, 16'hcdb5, 16'hcdb4, 16'hcd94, 16'hcd94, 16'hcd94, 16'hcd94, 16'hc594, 16'hc594, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc573, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb0, 16'h838c, 16'h3164, 16'h292, 16'h212, 16'h20e2, 16'h20e2, 16'h1081, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'ha4b1, 16'hacd2, 16'hacd2, 16'hb4d2, 16'hb4f2, 16'hb513, 16'hb513, 16'hb512, 16'hb512, 16'hb4f2, 16'hb512, 16'hb512, 16'had12, 16'hb532, 16'hb532, 16'hb553, 16'h9c90, 16'h5a89, 16'h8bee, 16'hacf2, 16'had12, 16'had12, 16'had12, 16'had12, 16'hacf2, 16'ha4d1, 16'h73b, 16'h6b2b, 16'h734c, 16'h62ca, 16'h8cf, 16'hbdb5, 16'ha4d2, 16'ha4b1, 16'h9c70, 16'h7b6b, 16'h7b4b, 16'h7b4b, 16'h838c, 16'h7b6b, 16'h20e2, 16'h841, 16'h841, 16'h18a2, 16'h1061, 16'h840, 16'h840, 16'h840, 16'h840, 16'h841, 16'h841, 16'h1041, 16'h4a28, 16'h83ee, 16'h5a68, 16'h527, 16'h5227, 16'h41a6, 16'h293, 16'h3144, 16'h41e7, 16'h5248, 16'h5228, 16'h5228, 16'h5227, 16'h4a8, 16'h4a7, 16'h4a27, 16'h4a7, 16'h49e7, 16'h49e7, 16'h49e6, 16'h49e6, 16'h49e6, 16'h39a5, 16'h20e3, 16'h1081, 16'h1061, 16'h840, 16'h840, 16'h840, 16'h840, 16'h840, 16'h020, 16'h020, 16'h020, 16'h18a1, 16'h3164, 16'h3143, 16'h3984, 16'h41a4, 16'h3984, 16'h3143, 16'h3964, 16'h41a4, 16'h3984, 16'h3984, 16'h3984, 16'h3984, 16'h3984, 16'h3984, 16'h3984, 16'h3984, 16'h3984, 16'h3984, 16'h3984, 16'h3984, 16'h3984, 16'h3184, 16'h3184, 16'h3984, 16'h3985, 16'h41a5, 16'h838d, 16'hee98, 16'heeb9, 16'heeb9, 16'heeb9, 16'heeb8, 16'he698, 16'he698, 16'he698, 16'he678, 16'he678, 16'hde77, 16'hde57, 16'hde57, 16'hde57, 16'hde57, 16'hde57, 16'hde57, 16'hde36, 16'hde16, 16'hde16, 16'hd616, 16'hd616, 16'hd5f6, 16'hd5f6, 16'hd5f6, 16'hd5f5, 16'hd5d5, 16'hcdd5, 16'hcdd5, 16'hcdb5, 16'hcdb5, 16'hcdb5, 16'hcdb4, 16'hcd94, 16'hcd94, 16'hc594, 16'hc594, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc573, 16'hc573, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4d2, 16'hb4d2, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'h83ad, 16'h3964, 16'h292, 16'h212, 16'h20e2, 16'h20e2, 16'h1081, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'ha470, 16'ha4b1, 16'hacb1, 16'hacb1, 16'hb4b2, 16'hb4f2, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb512, 16'hb532, 16'hb532, 16'hb533, 16'hb553, 16'h9c90, 16'h5a89, 16'h8ce, 16'had12, 16'hb533, 16'hb512, 16'had12, 16'had12, 16'had12, 16'hacf2, 16'h734c, 16'h4a7, 16'h5aca, 16'h39c6, 16'h5269, 16'h9450, 16'h9470, 16'h942f, 16'h8bee, 16'h7b4b, 16'h7b4b, 16'h7b4b, 16'h838c, 16'h7b6b, 16'h20c2, 16'h841, 16'h1061, 16'h5a89, 16'h5247, 16'h18a2, 16'h1081, 16'h1061, 16'h1081, 16'h1082, 16'h1882, 16'h18a2, 16'h213, 16'h3185, 16'h2924, 16'h294, 16'h49e6, 16'h5a68, 16'h6289, 16'h49e7, 16'h3124, 16'h41a6, 16'h5248, 16'h5a68, 16'h5248, 16'h5228, 16'h5228, 16'h5227, 16'h5227, 16'h4a28, 16'h5227, 16'h4a27, 16'h4a27, 16'h41c6, 16'h18c2, 16'h820, 16'h820, 16'h840, 16'h840, 16'h861, 16'h1081, 16'h10a2, 16'h18a2, 16'h10a1, 16'h1061, 16'h840, 16'h213, 16'h41c5, 16'h41a5, 16'h41a5, 16'h41a4, 16'h41a4, 16'h41a4, 16'h39a4, 16'h41a5, 16'h41e6, 16'h41e7, 16'h41e7, 16'h39c6, 16'h31a6, 16'h31a7, 16'h39c7, 16'h4a28, 16'h5248, 16'h4a48, 16'h4a48, 16'h5248, 16'h5269, 16'h5a89, 16'h5a89, 16'h5a89, 16'h5a89, 16'h5aaa, 16'h94f, 16'hee98, 16'heeb9, 16'heeb9, 16'heeb8, 16'he698, 16'he698, 16'he698, 16'he698, 16'he678, 16'hde77, 16'hde57, 16'hde57, 16'hde57, 16'hde37, 16'hde36, 16'hde37, 16'hde37, 16'hde36, 16'hd616, 16'hd616, 16'hd616, 16'hd5f6, 16'hd5f6, 16'hd5f6, 16'hd5f6, 16'hd5d5, 16'hd5d5, 16'hcdd5, 16'hcdb5, 16'hcdb5, 16'hcdb5, 16'hcdb4, 16'hcdb4, 16'hcd94, 16'hcd94, 16'hcd94, 16'hc594, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc553, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f2, 16'hb4d2, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'h83ad, 16'h3964, 16'h212, 16'h20e2, 16'h20e2, 16'h20e2, 16'h1081, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h9cf, 16'ha470, 16'ha4b1, 16'hacb1, 16'hacb1, 16'hacf2, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb512, 16'hb4f2, 16'hbd12, 16'hb553, 16'hb553, 16'hb553, 16'hbd73, 16'ha4b1, 16'h5a89, 16'h8ce, 16'hacd2, 16'hacf2, 16'ha4d1, 16'ha4b1, 16'h9c90, 16'h9c70, 16'h944f, 16'h734c, 16'h39c6, 16'h39e7, 16'h18e3, 16'h861, 16'h20e4, 16'h2924, 16'h294, 16'h41a6, 16'h73a, 16'h7b2b, 16'h7b4b, 16'h838c, 16'h736b, 16'h20c2, 16'h841, 16'h1061, 16'h7b6c, 16'h9c6f, 16'h5268, 16'h20e3, 16'h20c3, 16'h20e3, 16'h213, 16'h213, 16'h214, 16'h213, 16'h213, 16'h294, 16'h2924, 16'h6aea, 16'h8b6d, 16'hac91, 16'hac50, 16'h83b, 16'h49c6, 16'h3964, 16'h5248, 16'h5a68, 16'h62a9, 16'h6289, 16'h5248, 16'h5248, 16'h5248, 16'h5227, 16'h4a7, 16'h41c6, 16'h294, 16'h841, 16'h820, 16'h1061, 16'h18a2, 16'h20e2, 16'h213, 16'h213, 16'h2923, 16'h213, 16'h213, 16'h20e2, 16'h18a2, 16'h3144, 16'h49e5, 16'h41c5, 16'h41c5, 16'h41a5, 16'h41a4, 16'h41a4, 16'h41a5, 16'h41c5, 16'h5aa9, 16'h62ca, 16'h5aaa, 16'h52aa, 16'h4a8a, 16'h4a6a, 16'h526a, 16'h62ea, 16'h62ea, 16'h62ca, 16'h5aaa, 16'h62aa, 16'h62ca, 16'h62ca, 16'h62ea, 16'h62eb, 16'h62ca, 16'h62ea, 16'h942f, 16'hee98, 16'heeb9, 16'he698, 16'he698, 16'he698, 16'he698, 16'he698, 16'he678, 16'hde78, 16'hde77, 16'hde57, 16'hde57, 16'hde57, 16'hde37, 16'hde36, 16'hde36, 16'hde36, 16'hde36, 16'hd616, 16'hd616, 16'hd616, 16'hd5f6, 16'hd5f6, 16'hd5f5, 16'hd5f5, 16'hd5d5, 16'hcdd5, 16'hcdd5, 16'hcdd5, 16'hcdb5, 16'hcdb5, 16'hcdb4, 16'hcd94, 16'hcd94, 16'hc594, 16'hcd94, 16'hc594, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4d2, 16'hb4d2, 16'hb4d2, 16'hb4d1, 16'hb4d2, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacb1, 16'h8bad, 16'h3164, 16'h212, 16'h20e2, 16'h20e2, 16'h20e2, 16'h1081, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h93ce, 16'h9bef, 16'ha450, 16'ha4b1, 16'hacb1, 16'hacf2, 16'hb4f2, 16'hb4d2, 16'hb512, 16'hb4f2, 16'hbcd2, 16'hbd12, 16'hbd53, 16'hbd53, 16'hbd53, 16'hc594, 16'hacd1, 16'h5a89, 16'h6aeb, 16'h41e7, 16'h39a6, 16'h3185, 16'h3145, 16'h2924, 16'h214, 16'h213, 16'h18c3, 16'h18e3, 16'h2124, 16'h18c3, 16'h861, 16'h861, 16'h841, 16'h841, 16'h3124, 16'h73a, 16'h7b2b, 16'h7b4b, 16'h838c, 16'h7b6b, 16'h20c2, 16'h841, 16'h1061, 16'h7b6c, 16'hb532, 16'h83ee, 16'h5aa9, 16'h3144, 16'h20c3, 16'h18c2, 16'h18a2, 16'h18a2, 16'h18a2, 16'h18c2, 16'h18c2, 16'h20e3, 16'h6289, 16'h834c, 16'ha470, 16'hbc50, 16'hbc10, 16'h93ae, 16'h3124, 16'h3144, 16'h49e6, 16'h5248, 16'h6289, 16'h6289, 16'h5a69, 16'h5a68, 16'h5248, 16'h3164, 16'h2923, 16'h20e2, 16'h840, 16'h861, 16'h20e3, 16'h2923, 16'h2924, 16'h2924, 16'h2924, 16'h2923, 16'h2923, 16'h2923, 16'h293, 16'h293, 16'h3984, 16'h49c5, 16'h41a5, 16'h41c5, 16'h41c5, 16'h3984, 16'h3984, 16'h39a4, 16'h41c5, 16'h5aa9, 16'h5aca, 16'h5aaa, 16'h52aa, 16'h4a6a, 16'h4a6a, 16'h526a, 16'h62ca, 16'h62ca, 16'h5aaa, 16'h5aaa, 16'h5aaa, 16'h5aaa, 16'h62ca, 16'h62ea, 16'h62ca, 16'h62ca, 16'h62ca, 16'h942f, 16'he698, 16'heeb9, 16'he698, 16'he698, 16'he678, 16'he678, 16'hde78, 16'hde78, 16'hde57, 16'hde57, 16'hde57, 16'hde57, 16'hde57, 16'hde36, 16'hd636, 16'hd636, 16'hde36, 16'hd616, 16'hd616, 16'hd616, 16'hd5f6, 16'hd5f6, 16'hd5f6, 16'hd5d5, 16'hd5d5, 16'hcdd5, 16'hcdb5, 16'hcdb5, 16'hcdb5, 16'hcdb5, 16'hcd94, 16'hcd94, 16'hcd94, 16'hcd94, 16'hc594, 16'hc594, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc573, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4d2, 16'hb4d2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4d2, 16'hacd1, 16'h8bad, 16'h3964, 16'h213, 16'h20e2, 16'h20e2, 16'h20e2, 16'h1081, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h93ee, 16'h9ce, 16'h9c4f, 16'ha4b1, 16'hacb1, 16'hacd2, 16'hb4f2, 16'hb4f2, 16'hb4d2, 16'hbcf2, 16'hbd12, 16'hbd12, 16'hbd53, 16'hbd53, 16'hbd73, 16'hc594, 16'hacd1, 16'h5a89, 16'h62c9, 16'h18c2, 16'h1081, 16'h1061, 16'h1061, 16'h1061, 16'h1061, 16'h861, 16'h861, 16'h1082, 16'h213, 16'h18a2, 16'h840, 16'h841, 16'h1061, 16'h1062, 16'h3987, 16'h732b, 16'h7b2b, 16'h7b4b, 16'h838c, 16'h734a, 16'h213, 16'h1082, 16'h20e3, 16'h7b4c, 16'h9c90, 16'h83ae, 16'h8ce, 16'h5a88, 16'h213, 16'h18a2, 16'h18a2, 16'h18a2, 16'h18a3, 16'h18c3, 16'h20e3, 16'h20e3, 16'h5228, 16'h8bad, 16'ha42f, 16'hc451, 16'hcc11, 16'hb451, 16'h4a7, 16'h18a2, 16'h3124, 16'h3164, 16'h4a6, 16'h5a48, 16'h41a6, 16'h41c6, 16'h5268, 16'h213, 16'h18a2, 16'h861, 16'h820, 16'h18a2, 16'h2924, 16'h2923, 16'h3124, 16'h3144, 16'h3985, 16'h49e6, 16'h5247, 16'h62a9, 16'h62a9, 16'h6aea, 16'h6aea, 16'h49e6, 16'h41a5, 16'h41a4, 16'h41c5, 16'h3984, 16'h3964, 16'h39a4, 16'h41c5, 16'h5289, 16'h62ca, 16'h5aca, 16'h52aa, 16'h4a6a, 16'h4a6b, 16'h528a, 16'h62ca, 16'h5aaa, 16'h5aaa, 16'h5aaa, 16'h5aaa, 16'h5aaa, 16'h62ca, 16'h62ca, 16'h62ca, 16'h62ca, 16'h62ca, 16'h94f, 16'he678, 16'he698, 16'he698, 16'he678, 16'hde78, 16'hde78, 16'hde77, 16'hde57, 16'hde57, 16'hde57, 16'hde57, 16'hde37, 16'hde36, 16'hde36, 16'hd636, 16'hd616, 16'hd616, 16'hd616, 16'hd616, 16'hd616, 16'hd5f6, 16'hd5f5, 16'hd5d5, 16'hd5d5, 16'hd5d5, 16'hcdd5, 16'hcdb5, 16'hcdb5, 16'hcdb5, 16'hcdb4, 16'hcdb4, 16'hcd94, 16'hcd94, 16'hc594, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc573, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4d2, 16'hacd1, 16'h8bad, 16'h3964, 16'h212, 16'h20e2, 16'h20e2, 16'h20e2, 16'h1081, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h93cd, 16'h93ee, 16'h9ce, 16'ha470, 16'ha491, 16'hacb1, 16'hacd1, 16'hb512, 16'hb512, 16'hbcf2, 16'hbd33, 16'hbd53, 16'hc573, 16'hc573, 16'hc573, 16'hc594, 16'hacd1, 16'h6289, 16'h62c9, 16'h18e3, 16'h1061, 16'h1061, 16'h1061, 16'h1061, 16'h861, 16'h861, 16'h841, 16'h861, 16'h20e2, 16'h10a1, 16'h2924, 16'h49e6, 16'h527, 16'h3988, 16'h522b, 16'h6aea, 16'h73a, 16'h732a, 16'h7b4b, 16'h6ac9, 16'h3164, 16'h5247, 16'h5a88, 16'h6aca, 16'h6ac9, 16'h6aea, 16'h838c, 16'h838b, 16'h41c5, 16'h3984, 16'h41c5, 16'h41e6, 16'h41e6, 16'h49e6, 16'h49e6, 16'h49e6, 16'h527, 16'h93ce, 16'ha3ef, 16'hcc92, 16'hcc51, 16'hccb2, 16'h838d, 16'h41a6, 16'h20e3, 16'h20c2, 16'h39a5, 16'h5228, 16'h3164, 16'h3164, 16'h5268, 16'h3164, 16'h213, 16'h840, 16'h840, 16'h293, 16'h39a5, 16'h49c6, 16'h5a68, 16'h6aea, 16'h836c, 16'h8bcd, 16'h9c2e, 16'ha46f, 16'h9c2e, 16'h9c2f, 16'h8bcd, 16'h49e5, 16'h39a4, 16'h39a4, 16'h39a4, 16'h39a4, 16'h3984, 16'h41a4, 16'h3985, 16'h4a7, 16'h5aaa, 16'h5aca, 16'h528a, 16'h4a6a, 16'h528b, 16'h52ab, 16'h5aca, 16'h5aaa, 16'h5aaa, 16'h5aaa, 16'h5aaa, 16'h5aaa, 16'h5aaa, 16'h62ca, 16'h62ca, 16'h5aaa, 16'h62ca, 16'h942f, 16'hde57, 16'he678, 16'hde77, 16'hde77, 16'hde77, 16'hde57, 16'hde57, 16'hde57, 16'hde37, 16'hde37, 16'hde37, 16'hde36, 16'hde36, 16'hde36, 16'hd616, 16'hd616, 16'hd616, 16'hd5f6, 16'hd5f6, 16'hd5f6, 16'hd5f6, 16'hd5d5, 16'hd5d5, 16'hd5d5, 16'hcdd5, 16'hcdd5, 16'hcdb5, 16'hcdb5, 16'hcdb4, 16'hcd94, 16'hcd94, 16'hcd94, 16'hc594, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc573, 16'hc573, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4d2, 16'hacd1, 16'h8bcd, 16'h3964, 16'h292, 16'h20e2, 16'h20e2, 16'h20e2, 16'h1081, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h93cd, 16'h93ee, 16'h9c2f, 16'ha470, 16'hacb1, 16'hacb1, 16'hb4d2, 16'hb532, 16'hbd53, 16'hbd53, 16'hbd54, 16'hc553, 16'hc574, 16'hc574, 16'hc574, 16'hcdb4, 16'hacd1, 16'h6289, 16'h62c9, 16'h20e3, 16'h1061, 16'h1061, 16'h1061, 16'h1061, 16'h861, 16'h861, 16'h841, 16'h860, 16'h18c1, 16'h20e2, 16'h4a27, 16'h732a, 16'h6aca, 16'h4a2a, 16'h4ab, 16'h62aa, 16'h6ac9, 16'h732a, 16'h7b2a, 16'h6ac9, 16'h3964, 16'h6268, 16'h7b2a, 16'h7b2a, 16'h7b2b, 16'h7b2b, 16'h7b4b, 16'h7b6b, 16'h3984, 16'h20c2, 16'h20c2, 16'h20c2, 16'h18a2, 16'h18a2, 16'h1881, 16'h1881, 16'h20c3, 16'h838d, 16'hac30, 16'hdd97, 16'hdcd4, 16'hcc71, 16'hac50, 16'h8bad, 16'h5a89, 16'h3164, 16'h3985, 16'h41c6, 16'h2924, 16'h3164, 16'h5248, 16'h4a27, 16'h39e7, 16'h861, 16'h1061, 16'h4a7, 16'h73b, 16'h834c, 16'h93cd, 16'h94e, 16'h94e, 16'h93ee, 16'h93ed, 16'h93ee, 16'h8bcd, 16'h8bad, 16'h834b, 16'h49c5, 16'h3984, 16'h3984, 16'h3984, 16'h39a4, 16'h41a4, 16'h41a4, 16'h41a5, 16'h4a6, 16'h5a89, 16'h5aaa, 16'h528a, 16'h4a6a, 16'h4a8a, 16'h52ab, 16'h5aaa, 16'h5aaa, 16'h5aaa, 16'h5aaa, 16'h5aaa, 16'h5aaa, 16'h5aaa, 16'h5aaa, 16'h5aaa, 16'h5aaa, 16'h62ca, 16'h94f, 16'hde57, 16'hde77, 16'hde77, 16'hde57, 16'hde57, 16'hde57, 16'hde57, 16'hde37, 16'hde36, 16'hd636, 16'hd636, 16'hd616, 16'hd616, 16'hd616, 16'hd616, 16'hd5f6, 16'hd5f6, 16'hd5f6, 16'hd5f5, 16'hd5f5, 16'hd5d5, 16'hd5d5, 16'hd5d5, 16'hcdb5, 16'hcdb5, 16'hcdb5, 16'hcdb4, 16'hcdb4, 16'hcd94, 16'hcd94, 16'hcd94, 16'hc594, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc573, 16'hc573, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hacd2, 16'h8bcd, 16'h3984, 16'h292, 16'h20e2, 16'h20e2, 16'h20e2, 16'h1081, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h93ed, 16'h9bee, 16'h9c2f, 16'ha470, 16'hac91, 16'hac91, 16'hb4d2, 16'hb532, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hc573, 16'hc573, 16'hc574, 16'hcdb4, 16'hacf1, 16'h62a9, 16'h62c9, 16'h20e3, 16'h1061, 16'h1061, 16'h1061, 16'h1081, 16'h1061, 16'h861, 16'h861, 16'h861, 16'h18a1, 16'h20e2, 16'h41a6, 16'h5a68, 16'h49a5, 16'h28e4, 16'h3966, 16'h6aca, 16'h6aea, 16'h6288, 16'h6ae9, 16'h6b9, 16'h3144, 16'h49c6, 16'h7b2b, 16'h7b2b, 16'h7b2b, 16'h7b2b, 16'h7b4b, 16'h7b4b, 16'h3164, 16'h841, 16'h841, 16'h840, 16'h840, 16'h840, 16'h840, 16'h841, 16'h1862, 16'h72eb, 16'hc4d3, 16'he5f8, 16'hd4b3, 16'hc3f0, 16'hb471, 16'h8bad, 16'h6aca, 16'h41a5, 16'h3985, 16'h3965, 16'h294, 16'h3144, 16'h2944, 16'h39c6, 16'h5aaa, 16'h1061, 16'h1061, 16'h5a48, 16'h6aa9, 16'h834b, 16'h8bad, 16'h8bcd, 16'h8b8d, 16'h7b2b, 16'h73a, 16'h836c, 16'h7b4b, 16'h7b4b, 16'h73a, 16'h49c5, 16'h3984, 16'h3984, 16'h3984, 16'h3984, 16'h3984, 16'h39a4, 16'h39a4, 16'h4a6, 16'h5268, 16'h5a89, 16'h5269, 16'h4a6a, 16'h4a6a, 16'h526a, 16'h5aaa, 16'h5aaa, 16'h5aaa, 16'h5aaa, 16'h5aaa, 16'h5aaa, 16'h5aaa, 16'h5aaa, 16'h5aca, 16'h62aa, 16'h62ca, 16'h8cf, 16'hde37, 16'hde57, 16'hde57, 16'hde57, 16'hde37, 16'hde36, 16'hde36, 16'hde36, 16'hd616, 16'hd616, 16'hd616, 16'hd616, 16'hd616, 16'hd616, 16'hd5f6, 16'hd5f5, 16'hd5f5, 16'hd5d5, 16'hd5d5, 16'hd5d5, 16'hd5d5, 16'hd5d5, 16'hcdb5, 16'hcdb5, 16'hcdb5, 16'hcdb5, 16'hcdb4, 16'hcd94, 16'hcd94, 16'hcd94, 16'hc594, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc573, 16'hc573, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'h8bee, 16'h3984, 16'h292, 16'h212, 16'h20e2, 16'h20e2, 16'h1081, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h942e, 16'h9c2f, 16'ha42f, 16'hac70, 16'hac90, 16'hac71, 16'hb4f2, 16'hb512, 16'hbd32, 16'hbd53, 16'hbd53, 16'hbd32, 16'hbd73, 16'hbd73, 16'hc573, 16'hc5b4, 16'hacf1, 16'h6289, 16'h62c9, 16'h213, 16'h18c2, 16'h10a2, 16'h1081, 16'h1081, 16'h1081, 16'h1061, 16'h861, 16'h1081, 16'h861, 16'h1061, 16'h1081, 16'h1081, 16'h1061, 16'h1061, 16'h3144, 16'h73a, 16'h73b, 16'h49c6, 16'h732a, 16'h7b4a, 16'h20c2, 16'h49c6, 16'h7b2b, 16'h7b2b, 16'h7b2b, 16'h7b2b, 16'h7b4b, 16'h7b4a, 16'h3164, 16'h841, 16'h841, 16'h840, 16'h820, 16'h840, 16'h841, 16'h821, 16'h1842, 16'h7aab, 16'hd4f3, 16'hdcf4, 16'hcc31, 16'hc3cf, 16'hbc91, 16'h8bad, 16'h6aca, 16'h3985, 16'h3985, 16'h3965, 16'h293, 16'h3165, 16'h213, 16'h41c6, 16'h7b4c, 16'h18a2, 16'h1061, 16'h49c7, 16'h5a48, 16'h73a, 16'h7b2b, 16'h7b2b, 16'h73a, 16'h6289, 16'h5228, 16'h6aea, 16'h73a, 16'h72ea, 16'h6aca, 16'h49c5, 16'h3984, 16'h3984, 16'h3964, 16'h3984, 16'h3984, 16'h39a4, 16'h39a4, 16'h41c6, 16'h5227, 16'h5248, 16'h4a48, 16'h4a29, 16'h4a69, 16'h5a8a, 16'h5aaa, 16'h5a8a, 16'h5aaa, 16'h5aaa, 16'h5a8a, 16'h528a, 16'h5aaa, 16'h5aaa, 16'h62aa, 16'h62aa, 16'h62cb, 16'h8bef, 16'hd616, 16'hde37, 16'hde36, 16'hd636, 16'hd636, 16'hd616, 16'hd616, 16'hd616, 16'hd616, 16'hd616, 16'hd5f6, 16'hd5f6, 16'hd5f6, 16'hd5f6, 16'hd5d5, 16'hd5d5, 16'hd5d5, 16'hd5d5, 16'hd5d5, 16'hcdd5, 16'hcdd5, 16'hcdd5, 16'hcdb5, 16'hcdb5, 16'hcdb4, 16'hcd94, 16'hcd94, 16'hc594, 16'hc594, 16'hc594, 16'hc574, 16'hc574, 16'hc574, 16'hc573, 16'hc573, 16'hc573, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'h94e, 16'h3984, 16'h212, 16'h212, 16'h20e2, 16'h20e2, 16'h10a1, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h9c6f, 16'ha470, 16'hac70, 16'hacd1, 16'hb4f2, 16'hb4f2, 16'hb532, 16'hb532, 16'hbd32, 16'hbd53, 16'hbd53, 16'hbd12, 16'hbd53, 16'hc573, 16'hc573, 16'hc594, 16'hacf1, 16'h6289, 16'h62c9, 16'h213, 16'h18c2, 16'h1081, 16'h861, 16'h861, 16'h861, 16'h861, 16'h861, 16'h861, 16'h1081, 16'h10a2, 16'h1081, 16'h10a2, 16'h18c3, 16'h213, 16'h3984, 16'h6288, 16'h6ac9, 16'h4a7, 16'h5247, 16'h5247, 16'h2923, 16'h5227, 16'h7b2a, 16'h7b2b, 16'h7b2a, 16'h7b2a, 16'h7b4b, 16'h7b4a, 16'h3164, 16'h840, 16'h841, 16'h840, 16'h820, 16'h840, 16'h1061, 16'h1041, 16'h30a3, 16'hab8e, 16'he513, 16'hdc92, 16'hcc10, 16'hd410, 16'hc4b1, 16'h93ee, 16'h7b4c, 16'h3964, 16'h3144, 16'h3985, 16'h2924, 16'h3164, 16'h20e2, 16'h3985, 16'h62ca, 16'h18a2, 16'h841, 16'h2944, 16'h41c7, 16'h6289, 16'h72ea, 16'h6aca, 16'h6289, 16'h4a27, 16'h41e7, 16'h62a9, 16'h6aca, 16'h6aea, 16'h6289, 16'h41a5, 16'h3984, 16'h3984, 16'h3964, 16'h3984, 16'h3984, 16'h3984, 16'h41a5, 16'h39a5, 16'h49e6, 16'h41e6, 16'h49e6, 16'h41c6, 16'h49e6, 16'h5a47, 16'h62a9, 16'h62a9, 16'h5a89, 16'h528a, 16'h528a, 16'h528a, 16'h5aaa, 16'h5aaa, 16'h5aaa, 16'h62aa, 16'h62cb, 16'h8bee, 16'hd5f6, 16'hd616, 16'hd616, 16'hd616, 16'hd616, 16'hd616, 16'hd616, 16'hd5f6, 16'hd5f6, 16'hd5f6, 16'hd5f5, 16'hd5f5, 16'hd5f5, 16'hd5d5, 16'hcdd5, 16'hcdd5, 16'hcdd5, 16'hcdd5, 16'hcdb5, 16'hcdb5, 16'hcdb5, 16'hcdb5, 16'hcdb4, 16'hcd94, 16'hcd94, 16'hcd94, 16'hc594, 16'hc594, 16'hc594, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc553, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hb512, 16'hbd32, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'h942f, 16'h3985, 16'h292, 16'h20e2, 16'h20e2, 16'h20e2, 16'h10a1, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'ha4b0, 16'hacd1, 16'hacd1, 16'hb4f2, 16'hb532, 16'hb532, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd12, 16'hbd33, 16'hbd53, 16'hbd53, 16'hc574, 16'hacd1, 16'h6289, 16'h62a9, 16'h213, 16'h18e2, 16'h1081, 16'h861, 16'h861, 16'h861, 16'h861, 16'h860, 16'h861, 16'h213, 16'h2143, 16'h18c2, 16'h214, 16'h2945, 16'h2124, 16'h3164, 16'h6288, 16'h5227, 16'h4a6, 16'h49e6, 16'h4a27, 16'h292, 16'h49a5, 16'h7b2a, 16'h732b, 16'h7b2b, 16'h7b2b, 16'h7b4b, 16'h7b4a, 16'h3964, 16'h840, 16'h840, 16'h840, 16'h840, 16'h1081, 16'h5248, 16'h49c6, 16'h59c7, 16'hc410, 16'hd471, 16'hd410, 16'hd3f0, 16'he492, 16'hccb2, 16'h9cf, 16'h83ad, 16'h41a5, 16'h3124, 16'h3144, 16'h2924, 16'h2944, 16'h20e3, 16'h3165, 16'h5aa9, 16'h1061, 16'h840, 16'h2924, 16'h41c6, 16'h5228, 16'h6289, 16'h5a47, 16'h4a7, 16'h49e6, 16'h41c6, 16'h4a27, 16'h49e6, 16'h4a7, 16'h49e6, 16'h41c5, 16'h3984, 16'h3984, 16'h3164, 16'h3984, 16'h3984, 16'h3984, 16'h41a5, 16'h39a5, 16'h41c5, 16'h41c5, 16'h41e5, 16'h41c5, 16'h41c6, 16'h41c6, 16'h4a6, 16'h5a47, 16'h6288, 16'h62a9, 16'h5a89, 16'h5a8a, 16'h5aaa, 16'h5aaa, 16'h5aaa, 16'h5aaa, 16'h62ca, 16'h8bee, 16'hd5f5, 16'hd616, 16'hd5f6, 16'hd5f6, 16'hd5f6, 16'hd5f6, 16'hd5f6, 16'hd5f5, 16'hd5d5, 16'hd5d5, 16'hcdd5, 16'hcdd5, 16'hcdd5, 16'hcdd5, 16'hcdb5, 16'hcdb5, 16'hcdb5, 16'hcdb5, 16'hcdb5, 16'hcdb4, 16'hcdb4, 16'hcd94, 16'hcd94, 16'hc594, 16'hc594, 16'hc594, 16'hc594, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc553, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'h9c50, 16'h41a5, 16'h292, 16'h20e2, 16'h20e2, 16'h20e2, 16'h18a1, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'hacd1, 16'hacf1, 16'hb512, 16'hb532, 16'hb552, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd12, 16'hb512, 16'hb532, 16'hb532, 16'hbd33, 16'ha4b0, 16'h73b, 16'h6aea, 16'h213, 16'h18e2, 16'h10a1, 16'h861, 16'h861, 16'h861, 16'h861, 16'h860, 16'h861, 16'h1081, 16'h1081, 16'h1081, 16'h1081, 16'h10a2, 16'h10a2, 16'h3144, 16'h5a68, 16'h41c6, 16'h41a6, 16'h5247, 16'h62e9, 16'h18c3, 16'h4185, 16'h7ba, 16'h7b2b, 16'h73b, 16'h7b2b, 16'h7b4b, 16'h7b4a, 16'h3164, 16'h840, 16'h840, 16'h840, 16'h841, 16'h18a2, 16'h7b6c, 16'h94e, 16'h9bae, 16'hc410, 16'hd411, 16'hdc93, 16'he4b3, 16'hecf3, 16'hccb2, 16'h9c2f, 16'h8bad, 16'h41c6, 16'h3144, 16'h3144, 16'h2923, 16'h2944, 16'h213, 16'h3985, 16'h734c, 16'h18a2, 16'h841, 16'h3164, 16'h3165, 16'h3145, 16'h3164, 16'h3123, 16'h3984, 16'h41c5, 16'h3965, 16'h3144, 16'h3143, 16'h3164, 16'h49e6, 16'h41c5, 16'h3984, 16'h3984, 16'h3164, 16'h3964, 16'h3964, 16'h3984, 16'h39a4, 16'h39c5, 16'h41c5, 16'h41c5, 16'h41c6, 16'h41c6, 16'h41c6, 16'h41c6, 16'h49e6, 16'h49e6, 16'h49e6, 16'h5227, 16'h5a68, 16'h6289, 16'h5a89, 16'h528a, 16'h5a8a, 16'h5aaa, 16'h62ca, 16'h8bce, 16'hcdd5, 16'hd5f6, 16'hd5f6, 16'hd5f5, 16'hd5f5, 16'hd5d5, 16'hd5d5, 16'hd5d5, 16'hcdd5, 16'hcdd5, 16'hcdd5, 16'hcdd5, 16'hcdb5, 16'hcdb5, 16'hcdb5, 16'hcdb5, 16'hcdb4, 16'hcd94, 16'hcd94, 16'hcd94, 16'hcd94, 16'hc594, 16'hc594, 16'hc594, 16'hc594, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc573, 16'hc573, 16'hc573, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'h9c50, 16'h4185, 16'h292, 16'h212, 16'h20e2, 16'h20e2, 16'h18a1, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'hacd1, 16'hacf1, 16'hacf2, 16'had12, 16'hb512, 16'hacf2, 16'hacf2, 16'hacd1, 16'hacd1, 16'ha4b1, 16'ha491, 16'ha490, 16'h9c70, 16'h9c70, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h944f, 16'h7b6c, 16'h213, 16'h20e3, 16'h10a2, 16'h861, 16'h861, 16'h861, 16'h861, 16'h861, 16'h861, 16'h10a1, 16'h10a1, 16'h10a1, 16'h10a1, 16'h18c2, 16'h18e2, 16'h3144, 16'h6ac9, 16'h5a68, 16'h41a6, 16'h5227, 16'h62cb, 16'h2948, 16'h49a8, 16'h7bb, 16'h7b2b, 16'h7bb, 16'h7bb, 16'h7b4b, 16'h7b4a, 16'h3164, 16'h820, 16'h840, 16'h841, 16'h1061, 16'h20a2, 16'h73a, 16'h9c2f, 16'hc512, 16'hc410, 16'hdc93, 16'hee5a, 16'hf5d7, 16'he513, 16'hc4b2, 16'ha450, 16'h8bad, 16'h41a5, 16'h3144, 16'h3164, 16'h2923, 16'h2924, 16'h2924, 16'h3985, 16'h732c, 16'h18c3, 16'h841, 16'h3164, 16'h2924, 16'h41c6, 16'h426, 16'h41c6, 16'h41e6, 16'h41a5, 16'h3985, 16'h41c6, 16'h4a7, 16'h5247, 16'h6288, 16'h49c5, 16'h3984, 16'h3983, 16'h3963, 16'h3964, 16'h3964, 16'h3984, 16'h39a4, 16'h3164, 16'h3124, 16'h3985, 16'h49c6, 16'h49e6, 16'h41c6, 16'h41c6, 16'h49c5, 16'h49e6, 16'h49e6, 16'h49e6, 16'h49e6, 16'h5226, 16'h5a67, 16'h5a89, 16'h5a69, 16'h5a89, 16'h62ca, 16'h8bce, 16'hcdb5, 16'hd5d5, 16'hd5d5, 16'hcdd5, 16'hcdd5, 16'hcdd5, 16'hcdd5, 16'hcdd5, 16'hcdd5, 16'hcdb5, 16'hcdb5, 16'hcdb5, 16'hcdb5, 16'hcdb4, 16'hcd94, 16'hcd94, 16'hcd94, 16'hcd94, 16'hc594, 16'hc594, 16'hc594, 16'hc594, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc573, 16'hc573, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb512, 16'hb512, 16'hb4f2, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'h9c30, 16'h3985, 16'h292, 16'h212, 16'h20e2, 16'h20e2, 16'h18a1, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'ha4b0, 16'ha4d1, 16'hacd1, 16'hacf1, 16'hacf1, 16'hacf2, 16'hacd2, 16'hacd1, 16'hacd1, 16'ha4b1, 16'ha4b1, 16'ha4b0, 16'ha490, 16'ha490, 16'h9c70, 16'h9c70, 16'h9c50, 16'h9c4f, 16'h7b6c, 16'h213, 16'h213, 16'h18a2, 16'h861, 16'h860, 16'h861, 16'h861, 16'h861, 16'h861, 16'h860, 16'h840, 16'h860, 16'h861, 16'h1061, 16'h1081, 16'h3124, 16'h6ae9, 16'h62a8, 16'h73a, 16'h7b4b, 16'h5269, 16'h2949, 16'h49c9, 16'h73b, 16'h73a, 16'h7ba, 16'h7b2a, 16'h7b4b, 16'h7b2a, 16'h3164, 16'h820, 16'h840, 16'h1041, 16'h1061, 16'h1882, 16'h836c, 16'ha42f, 16'hccf3, 16'hd492, 16'he4d4, 16'hf6db, 16'hf596, 16'hd4b2, 16'hc4d2, 16'ha470, 16'h8bce, 16'h49e6, 16'h2923, 16'h3143, 16'h2923, 16'h2924, 16'h2924, 16'h3185, 16'h62ca, 16'h18c2, 16'h861, 16'h3985, 16'h41a6, 16'h39a5, 16'h4a7, 16'h41c6, 16'h41c5, 16'h5227, 16'h5a68, 16'h5a88, 16'h6289, 16'h6289, 16'h62a9, 16'h49c5, 16'h3984, 16'h3983, 16'h3963, 16'h3984, 16'h3964, 16'h3984, 16'h3984, 16'h3164, 16'h2923, 16'h2923, 16'h3144, 16'h39a5, 16'h49c6, 16'h41c5, 16'h5246, 16'h5226, 16'h41c5, 16'h4185, 16'h4184, 16'h41a4, 16'h41a4, 16'h49c4, 16'h41a4, 16'h4a7, 16'h5aaa, 16'h83ce, 16'hcdb4, 16'hcdd5, 16'hcdd5, 16'hcdd5, 16'hcdb5, 16'hcdb5, 16'hcdb5, 16'hcdb5, 16'hcdb5, 16'hcdb5, 16'hcdb5, 16'hcdb4, 16'hcd94, 16'hcd94, 16'hc594, 16'hc594, 16'hc594, 16'hc594, 16'hc594, 16'hc594, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc573, 16'hc553, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hbd32, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'h9c50, 16'h41a5, 16'h212, 16'h212, 16'h20e2, 16'h20e2, 16'h18a1, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'ha490, 16'ha4b1, 16'ha4b1, 16'hacd1, 16'hacd1, 16'ha4b1, 16'ha4b1, 16'ha4b1, 16'ha4b1, 16'ha4b1, 16'ha4b0, 16'ha4b0, 16'ha4b0, 16'ha4b1, 16'ha4b1, 16'hacd1, 16'h9c50, 16'h73b, 16'h6aea, 16'h213, 16'h213, 16'h18a2, 16'h861, 16'h860, 16'h861, 16'h861, 16'h861, 16'h860, 16'h860, 16'h840, 16'h212, 16'h2123, 16'h840, 16'h861, 16'h3124, 16'h73a, 16'h6288, 16'h5a88, 16'h732b, 16'h732b, 16'h4ab, 16'h52b, 16'h73b, 16'h732a, 16'h7b2a, 16'h7b2a, 16'h7b4b, 16'h7b2a, 16'h3164, 16'h820, 16'h840, 16'h841, 16'h1061, 16'h20c3, 16'h83ad, 16'hb4d1, 16'hd554, 16'he514, 16'he4f4, 16'hf65a, 16'hed34, 16'hc470, 16'hc513, 16'h9c50, 16'h8bcd, 16'h5227, 16'h3144, 16'h2923, 16'h293, 16'h213, 16'h2924, 16'h3165, 16'h5a89, 16'h1082, 16'h840, 16'h3985, 16'h5247, 16'h5227, 16'h49c6, 16'h3985, 16'h3164, 16'h49e6, 16'h4a6, 16'h5247, 16'h5a68, 16'h5a69, 16'h6288, 16'h41c5, 16'h3984, 16'h3983, 16'h3983, 16'h3984, 16'h3964, 16'h3984, 16'h39a4, 16'h41c5, 16'h3164, 16'h3184, 16'h3985, 16'h3164, 16'h41a5, 16'h4a6, 16'h49e5, 16'h3122, 16'h312, 16'h312, 16'h312, 16'h311, 16'h30e1, 16'h30e1, 16'h311, 16'h3923, 16'h41e7, 16'h838d, 16'hc594, 16'hcdb5, 16'hcdb5, 16'hcdb5, 16'hcdb4, 16'hcdb5, 16'hcdb5, 16'hcdb5, 16'hcdb4, 16'hcd94, 16'hcd94, 16'hcd94, 16'hcd94, 16'hc594, 16'hc594, 16'hc594, 16'hc594, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc573, 16'hc573, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hbd33, 16'hbd33, 16'hbd33, 16'hb512, 16'hb512, 16'h9c70, 16'h41a5, 16'h213, 16'h212, 16'h20e2, 16'h20e2, 16'h18a1, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'hb532, 16'hb532, 16'hb532, 16'hb532, 16'hbd53, 16'hb553, 16'hb553, 16'hb533, 16'hb533, 16'hb533, 16'hb532, 16'had12, 16'had12, 16'hb512, 16'hb512, 16'hb533, 16'hacb1, 16'h62a9, 16'h62c9, 16'h213, 16'h213, 16'h18a2, 16'h1061, 16'h861, 16'h861, 16'h861, 16'h861, 16'h861, 16'h860, 16'h840, 16'h1081, 16'h1081, 16'h840, 16'h1081, 16'h3964, 16'h73a, 16'h732a, 16'h6aea, 16'h6aca, 16'h62a9, 16'h5a6b, 16'h5a4b, 16'h73a, 16'h732a, 16'h7ba, 16'h7b2a, 16'h7b4b, 16'h7b2a, 16'h3164, 16'h820, 16'h821, 16'h841, 16'h1882, 16'h49c7, 16'h93ee, 16'ha470, 16'hd555, 16'hdcd4, 16'hed56, 16'hf619, 16'he4d3, 16'hbc50, 16'hbd33, 16'h9c50, 16'h8bce, 16'h5247, 16'h3164, 16'h2923, 16'h213, 16'h20e3, 16'h213, 16'h3165, 16'h4a48, 16'h1082, 16'h840, 16'h3184, 16'h5227, 16'h4a7, 16'h3985, 16'h3164, 16'h3164, 16'h41c6, 16'h5227, 16'h5a48, 16'h5a68, 16'h5a68, 16'h5a88, 16'h41c5, 16'h3984, 16'h3984, 16'h3964, 16'h3163, 16'h3983, 16'h3984, 16'h49e6, 16'h5227, 16'h41a5, 16'h5226, 16'h5a67, 16'h6287, 16'h6aa7, 16'h5a67, 16'h3143, 16'h2081, 16'h28c1, 16'h28a1, 16'h28a1, 16'h20a1, 16'h20a0, 16'h20a1, 16'h28c1, 16'h20a1, 16'h3164, 16'h732c, 16'hc574, 16'hcdb5, 16'hcdb5, 16'hcd94, 16'hcd94, 16'hcd94, 16'hcd94, 16'hcd94, 16'hcd94, 16'hcd94, 16'hcd94, 16'hc594, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc573, 16'hc553, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hbd12, 16'hbd12, 16'hbd33, 16'hb513, 16'hb512, 16'hb512, 16'ha491, 16'h41a6, 16'h213, 16'h212, 16'h20e2, 16'h20e2, 16'h1881, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'hbd53, 16'hbd53, 16'had32, 16'had32, 16'hb553, 16'hbd53, 16'hb553, 16'hb533, 16'hb533, 16'hb533, 16'hb533, 16'had12, 16'had12, 16'hb512, 16'hb512, 16'hb533, 16'hacd1, 16'h62a9, 16'h62c9, 16'h213, 16'h213, 16'h18c2, 16'h1061, 16'h1061, 16'h861, 16'h861, 16'h861, 16'h860, 16'h860, 16'h840, 16'h840, 16'h020, 16'h840, 16'h10a2, 16'h3944, 16'h73a, 16'h7b2a, 16'h7b2a, 16'h7b6c, 16'h6289, 16'h41a6, 16'h5a48, 16'h73a, 16'h73a, 16'h73a, 16'h7b2a, 16'h7b4a, 16'h7b2a, 16'h3164, 16'h820, 16'h841, 16'h294, 16'h528, 16'h62a9, 16'h7b4c, 16'h832c, 16'hcc92, 16'hdc93, 16'hedf8, 16'hed96, 16'he4d3, 16'hb491, 16'hb4b1, 16'h9c50, 16'h8bcd, 16'h49e7, 16'h3144, 16'h3144, 16'h2923, 16'h18c2, 16'h213, 16'h3165, 16'h4a8, 16'h1081, 16'h840, 16'h3184, 16'h5227, 16'h5247, 16'h49e6, 16'h3985, 16'h49e6, 16'h5227, 16'h5a48, 16'h5247, 16'h5227, 16'h5248, 16'h5a68, 16'h41c5, 16'h3984, 16'h3984, 16'h3984, 16'h3143, 16'h3143, 16'h3164, 16'h3163, 16'h2943, 16'h293, 16'h293, 16'h313, 16'h5a46, 16'h6266, 16'h3984, 16'h1061, 16'h1060, 16'h20a1, 16'h20c1, 16'h20c1, 16'h20a1, 16'h1061, 16'h1061, 16'h1881, 16'h1881, 16'h2924, 16'h6aeb, 16'hc574, 16'hcd94, 16'hcd94, 16'hcd94, 16'hcd94, 16'hc574, 16'hc574, 16'hc594, 16'hc594, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc573, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hbd33, 16'hbd33, 16'hb512, 16'hb512, 16'ha4b1, 16'h41a6, 16'h293, 16'h212, 16'h20e2, 16'h20e2, 16'h18a1, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'hbd53, 16'hbd53, 16'hb532, 16'hb552, 16'hbd53, 16'hbd53, 16'hb533, 16'hb532, 16'had12, 16'had32, 16'hb533, 16'had12, 16'had12, 16'had12, 16'had12, 16'hb532, 16'hacd1, 16'h62a9, 16'h6aca, 16'h3985, 16'h3164, 16'h18c2, 16'h1081, 16'h1061, 16'h1061, 16'h861, 16'h861, 16'h860, 16'h840, 16'h840, 16'h840, 16'h840, 16'h840, 16'h1081, 16'h3144, 16'h72e9, 16'h739, 16'h6ae9, 16'h732a, 16'h6ac9, 16'h5a66, 16'h7b27, 16'h7ba, 16'h73a, 16'h73a, 16'h7b2a, 16'h7b2a, 16'h7b2a, 16'h3144, 16'h840, 16'h841, 16'h3125, 16'h7b2c, 16'h73a, 16'h6a88, 16'h7aea, 16'hccd2, 16'hdd14, 16'hee18, 16'hecf3, 16'hdcf3, 16'hbcb1, 16'hb4d2, 16'h9c4f, 16'h8bad, 16'h49c6, 16'h2923, 16'h3144, 16'h2924, 16'h18a2, 16'h20e3, 16'h3145, 16'h427, 16'h1061, 16'h840, 16'h3164, 16'h4a6, 16'h527, 16'h5227, 16'h5247, 16'h5a68, 16'h5a68, 16'h5a48, 16'h5a48, 16'h5227, 16'h5227, 16'h5a68, 16'h41c5, 16'h3984, 16'h3984, 16'h3984, 16'h3143, 16'h3163, 16'h3164, 16'h3143, 16'h20e2, 16'h18c2, 16'h1881, 16'h293, 16'h51e5, 16'h51e4, 16'h525, 16'h293, 16'h1061, 16'h292, 16'h292, 16'h20c2, 16'h20a2, 16'h18a1, 16'h1061, 16'h1061, 16'h1881, 16'h2924, 16'h6aea, 16'hc553, 16'hc594, 16'hc594, 16'hc594, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc573, 16'hc573, 16'hc573, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hbd32, 16'hbd33, 16'hbd33, 16'hb512, 16'hb512, 16'hacb1, 16'h41c6, 16'h293, 16'h212, 16'h20e2, 16'h20e2, 16'h18a1, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'hbd53, 16'hbd53, 16'hb552, 16'hb552, 16'hb553, 16'hbd53, 16'hb532, 16'had32, 16'had12, 16'hb532, 16'hb532, 16'had32, 16'ha512, 16'had12, 16'had12, 16'hb532, 16'hacb1, 16'h62a9, 16'h8bce, 16'h942f, 16'h5ac9, 16'h18e2, 16'h1081, 16'h1081, 16'h1081, 16'h1081, 16'h1081, 16'h1081, 16'h881, 16'h861, 16'h860, 16'h841, 16'h841, 16'h861, 16'h18a2, 16'h3144, 16'h2923, 16'h213, 16'h20e2, 16'h18c2, 16'h20c2, 16'h51e5, 16'h73a, 16'h73a, 16'h73a, 16'h7ba, 16'h7b2b, 16'h7b2a, 16'h3143, 16'h840, 16'h840, 16'h1061, 16'h41c6, 16'h7b2a, 16'h6aa8, 16'h83a, 16'hcc31, 16'he515, 16'hedb7, 16'he492, 16'he574, 16'hbcd2, 16'hbd33, 16'h9c2f, 16'h8bcd, 16'h5227, 16'h3124, 16'h2923, 16'h293, 16'h1081, 16'h18c2, 16'h2944, 16'h41e7, 16'h1061, 16'h840, 16'h3164, 16'h49e6, 16'h527, 16'h5227, 16'h5a48, 16'h5a47, 16'h5a47, 16'h5247, 16'h5227, 16'h527, 16'h5227, 16'h5a47, 16'h41c5, 16'h3984, 16'h3984, 16'h3964, 16'h3964, 16'h3164, 16'h3964, 16'h3163, 16'h293, 16'h1061, 16'h1881, 16'h3984, 16'h20e2, 16'h20c1, 16'h41c4, 16'h49e5, 16'h20e2, 16'h20e1, 16'h28e2, 16'h28e2, 16'h28e2, 16'h292, 16'h20e2, 16'h20c2, 16'h3123, 16'h3985, 16'h6aca, 16'hbd53, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc573, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hbd32, 16'hbd33, 16'hb532, 16'hbd32, 16'hb512, 16'hacf2, 16'h41c6, 16'h293, 16'h212, 16'h20e2, 16'h20e2, 16'h18a1, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'hbd52, 16'hb532, 16'hb532, 16'hb553, 16'hb553, 16'hbd53, 16'hb553, 16'hb532, 16'hb533, 16'hb533, 16'hb532, 16'had32, 16'ha512, 16'had12, 16'had12, 16'hb532, 16'ha4b1, 16'h62a9, 16'h94e, 16'ha4b0, 16'h62e9, 16'h18c2, 16'h1081, 16'h10a1, 16'h861, 16'h861, 16'h861, 16'h861, 16'h861, 16'h860, 16'h860, 16'h841, 16'h840, 16'h840, 16'h841, 16'h841, 16'h861, 16'h840, 16'h860, 16'h840, 16'h840, 16'h4165, 16'h72ea, 16'h73a, 16'h73a, 16'h73a, 16'h7b2b, 16'h732a, 16'h2943, 16'h840, 16'h841, 16'h1041, 16'h1882, 16'h6ac9, 16'h6aa8, 16'h8ba, 16'hbbcf, 16'he535, 16'hed96, 16'he4b2, 16'he595, 16'hb4b1, 16'hbd33, 16'h9c2f, 16'h8bce, 16'h5248, 16'h3164, 16'h2944, 16'h213, 16'h1061, 16'h18c2, 16'h2944, 16'h39a6, 16'h861, 16'h840, 16'h2943, 16'h41c5, 16'h49e5, 16'h49e5, 16'h41c5, 16'h49c5, 16'h526, 16'h41a5, 16'h3984, 16'h49e5, 16'h5227, 16'h6aa9, 16'h41a5, 16'h3984, 16'h3984, 16'h3964, 16'h3163, 16'h3163, 16'h3964, 16'h3143, 16'h2923, 16'h1081, 16'h293, 16'h3144, 16'h841, 16'h840, 16'h1081, 16'h3163, 16'h41a4, 16'h3123, 16'h3963, 16'h3963, 16'h3963, 16'h3963, 16'h3123, 16'h3122, 16'h3963, 16'h3985, 16'h6aca, 16'hbd53, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc574, 16'hc573, 16'hc573, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hb532, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hb513, 16'hb4f2, 16'h49c7, 16'h293, 16'h212, 16'h20e2, 16'h20e2, 16'h18a1, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'hb512, 16'hacd1, 16'hb532, 16'hbd53, 16'hbd53, 16'hbd53, 16'hb532, 16'hb512, 16'hb532, 16'hb533, 16'hb532, 16'had12, 16'h9d11, 16'had12, 16'had12, 16'hb532, 16'ha4b1, 16'h62a9, 16'h94e, 16'ha4b0, 16'h62c9, 16'h18c2, 16'h1081, 16'h18c2, 16'h1081, 16'h861, 16'h861, 16'h861, 16'h861, 16'h861, 16'h861, 16'h861, 16'h861, 16'h861, 16'h861, 16'h861, 16'h841, 16'h841, 16'h840, 16'h840, 16'h840, 16'h4185, 16'h72ea, 16'h73a, 16'h73a, 16'h73a, 16'h6ac9, 16'h5a48, 16'h3164, 16'h20e3, 16'h20e3, 16'h2924, 16'h41a4, 16'h7b9, 16'h72a9, 16'h932c, 16'hc410, 16'he535, 16'he4d3, 16'he4f3, 16'hdd95, 16'hb4b1, 16'hbd53, 16'h9c50, 16'h8bce, 16'h4a7, 16'h3144, 16'h3144, 16'h293, 16'h1081, 16'h18a2, 16'h2924, 16'h3185, 16'h861, 16'h820, 16'h292, 16'h3983, 16'h3983, 16'h2923, 16'h20e2, 16'h3123, 16'h49c5, 16'h3143, 16'h2923, 16'h49c6, 16'h5a28, 16'h72ea, 16'h41c5, 16'h3984, 16'h3984, 16'h3984, 16'h3183, 16'h3164, 16'h3163, 16'h3143, 16'h2923, 16'h20e2, 16'h3164, 16'h20c2, 16'h841, 16'h861, 16'h1061, 16'h18a1, 16'h41a4, 16'h41a4, 16'h3963, 16'h3963, 16'h3963, 16'h3943, 16'h3123, 16'h3122, 16'h3964, 16'h3985, 16'h62ca, 16'hbd53, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc573, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hb532, 16'hb532, 16'hb532, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hacd1, 16'hb4d1, 16'hb4d1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f2, 16'hb4f1, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hbd33, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'h49e7, 16'h293, 16'h212, 16'h20e2, 16'h20e2, 16'h18a1, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'hb532, 16'hacf1, 16'hb532, 16'hb512, 16'hb532, 16'hb512, 16'hb512, 16'hb512, 16'hb532, 16'hb533, 16'hb533, 16'had12, 16'ha512, 16'hb512, 16'hb512, 16'hb532, 16'ha4b0, 16'h62a9, 16'h8ce, 16'ha4b0, 16'h62c9, 16'h18c2, 16'h1081, 16'h20c2, 16'h10a1, 16'h861, 16'h861, 16'h861, 16'h861, 16'h861, 16'h861, 16'h861, 16'h861, 16'h861, 16'h861, 16'h841, 16'h840, 16'h840, 16'h840, 16'h840, 16'h840, 16'h4185, 16'h72ea, 16'h73a, 16'h73a, 16'h73a, 16'h7b2a, 16'h6ac9, 16'h3144, 16'h1081, 16'h20c3, 16'h3144, 16'h526, 16'h7b2a, 16'h6aa9, 16'h93c, 16'hc410, 16'hd472, 16'hcc10, 16'hdd13, 16'hddb5, 16'hbcf2, 16'hc554, 16'h9c50, 16'h93ce, 16'h5a48, 16'h2923, 16'h2923, 16'h2923, 16'h1081, 16'h18a2, 16'h213, 16'h3185, 16'h861, 16'h820, 16'h20e2, 16'h3143, 16'h3143, 16'h3143, 16'h2923, 16'h3143, 16'h3123, 16'h2923, 16'h3144, 16'h5227, 16'h6a89, 16'h72ea, 16'h41a5, 16'h3984, 16'h3984, 16'h3983, 16'h3183, 16'h3164, 16'h3164, 16'h3143, 16'h293, 16'h3144, 16'h2923, 16'h1061, 16'h840, 16'h861, 16'h840, 16'h1061, 16'h3123, 16'h5a46, 16'h49e4, 16'h4163, 16'h3963, 16'h3943, 16'h3143, 16'h3123, 16'h3964, 16'h3985, 16'h62aa, 16'hbd33, 16'hc553, 16'hc553, 16'hc573, 16'hc573, 16'hc573, 16'hc553, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hacd1, 16'hb4d1, 16'hb4d1, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hbd32, 16'hb512, 16'hb512, 16'hb512, 16'hbd13, 16'hb513, 16'h49e7, 16'h293, 16'h213, 16'h20e2, 16'h20e2, 16'h18a1, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'hbd53, 16'hbd33, 16'hbd53, 16'hb512, 16'hb512, 16'hacf2, 16'hb512, 16'hb512, 16'hb532, 16'hb533, 16'hb533, 16'had32, 16'had32, 16'hb532, 16'hb532, 16'hb532, 16'ha490, 16'h62a9, 16'h94e, 16'ha490, 16'h62c9, 16'h18c2, 16'h1081, 16'h20c2, 16'h10a2, 16'h840, 16'h860, 16'h861, 16'h861, 16'h861, 16'h861, 16'h861, 16'h861, 16'h841, 16'h840, 16'h840, 16'h020, 16'h820, 16'h840, 16'h841, 16'h841, 16'h4185, 16'h72e9, 16'h72ea, 16'h72ea, 16'h73a, 16'h7b2a, 16'h739, 16'h2923, 16'h820, 16'h820, 16'h840, 16'h20a2, 16'h6aa8, 16'h6aa9, 16'h82ca, 16'hc3ef, 16'hbbaf, 16'h9bc, 16'hccd2, 16'hddb5, 16'hb4d2, 16'hbd53, 16'h9c50, 16'h8bad, 16'h5a48, 16'h3164, 16'h2923, 16'h213, 16'h1081, 16'h18a2, 16'h18e3, 16'h2965, 16'h861, 16'h820, 16'h1081, 16'h18c2, 16'h18a1, 16'h18c2, 16'h20e2, 16'h293, 16'h2923, 16'h2923, 16'h3164, 16'h5247, 16'h6a89, 16'h73a, 16'h41c5, 16'h3984, 16'h3983, 16'h3983, 16'h3183, 16'h3163, 16'h3164, 16'h3143, 16'h2923, 16'h3164, 16'h18a2, 16'h820, 16'h820, 16'h820, 16'h820, 16'h840, 16'h20c2, 16'h49c4, 16'h5a46, 16'h49e5, 16'h4163, 16'h3943, 16'h3143, 16'h3123, 16'h3964, 16'h3985, 16'h62aa, 16'hbd32, 16'hc553, 16'hc553, 16'hc553, 16'hc553, 16'hc553, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d2, 16'hb4d1, 16'hb4d1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb513, 16'hb4f3, 16'h49e7, 16'h293, 16'h213, 16'h20e2, 16'h20e2, 16'h18a1, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'hbd53, 16'hbd53, 16'hbd52, 16'hb532, 16'hb532, 16'hb512, 16'hb512, 16'hacf1, 16'hb512, 16'hb533, 16'hb532, 16'had12, 16'had12, 16'hb532, 16'hb532, 16'hb532, 16'h9c8f, 16'h62a9, 16'h94e, 16'h9c90, 16'h62c9, 16'h18a2, 16'h1081, 16'h20e2, 16'h18c2, 16'h840, 16'h840, 16'h860, 16'h860, 16'h861, 16'h860, 16'h860, 16'h840, 16'h840, 16'h840, 16'h840, 16'h840, 16'h841, 16'h861, 16'h10a1, 16'h861, 16'h3984, 16'h72e9, 16'h72ea, 16'h72ea, 16'h72e9, 16'h7b2a, 16'h739, 16'h2923, 16'h840, 16'h840, 16'h840, 16'h1861, 16'h6268, 16'h6aa9, 16'h7aca, 16'hbce, 16'habce, 16'h82eb, 16'hb450, 16'hd5b5, 16'hacb1, 16'hbd53, 16'h9c30, 16'h8bad, 16'h5227, 16'h3964, 16'h3144, 16'h213, 16'h1061, 16'h1081, 16'h18c2, 16'h2924, 16'h841, 16'h820, 16'h20e2, 16'h3963, 16'h3984, 16'h3984, 16'h3963, 16'h3143, 16'h2922, 16'h20e2, 16'h2923, 16'h5227, 16'h6a89, 16'h73b, 16'h41c5, 16'h3984, 16'h3983, 16'h3964, 16'h3163, 16'h3163, 16'h3163, 16'h3163, 16'h2943, 16'h213, 16'h840, 16'h820, 16'h820, 16'h820, 16'h820, 16'h840, 16'h20e1, 16'h3963, 16'h49e4, 16'h525, 16'h41a4, 16'h3963, 16'h3943, 16'h3143, 16'h3964, 16'h3965, 16'h62a9, 16'hbd32, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hb4d1, 16'hb4f1, 16'hb4d1, 16'hb4f1, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb532, 16'hb512, 16'hb4f2, 16'h49e7, 16'h293, 16'h213, 16'h20e2, 16'h20e2, 16'h18a1, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'hbd53, 16'hb533, 16'hb532, 16'hb532, 16'hb512, 16'hacf2, 16'hacd1, 16'hacd1, 16'hb4f2, 16'hb532, 16'hb532, 16'had12, 16'had12, 16'hb532, 16'hb532, 16'hb532, 16'h9c6f, 16'h62a9, 16'h942e, 16'h9c90, 16'h62ea, 16'h18a2, 16'h1081, 16'h20e3, 16'h18c2, 16'h840, 16'h840, 16'h840, 16'h861, 16'h841, 16'h861, 16'h860, 16'h840, 16'h840, 16'h840, 16'h840, 16'h840, 16'h861, 16'h1061, 16'h20e3, 16'h1061, 16'h3984, 16'h6ae9, 16'h72e9, 16'h72e9, 16'h72ea, 16'h7b2a, 16'h739, 16'h2923, 16'h820, 16'h841, 16'h1882, 16'h20c2, 16'h6288, 16'h6aa9, 16'h72ca, 16'h9bad, 16'hac2f, 16'h93ce, 16'ha4f, 16'hc553, 16'hac91, 16'hbd53, 16'h9cf, 16'h838d, 16'h49c6, 16'h3123, 16'h3144, 16'h2924, 16'h1081, 16'h1081, 16'h18a2, 16'h213, 16'h841, 16'h820, 16'h20e2, 16'h3963, 16'h4184, 16'h4184, 16'h3984, 16'h3964, 16'h3143, 16'h3143, 16'h3164, 16'h5227, 16'h6aa9, 16'h73b, 16'h41a4, 16'h3984, 16'h3984, 16'h3984, 16'h3143, 16'h3143, 16'h3163, 16'h3984, 16'h20e2, 16'h861, 16'h820, 16'h820, 16'h820, 16'h820, 16'h820, 16'h840, 16'h20c2, 16'h3943, 16'h3943, 16'h3963, 16'h3963, 16'h3942, 16'h3943, 16'h3142, 16'h3964, 16'h3985, 16'h62a9, 16'hbd32, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hb4d1, 16'hb4d1, 16'hb4d2, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb513, 16'h4a7, 16'h293, 16'h293, 16'h20e2, 16'h20e2, 16'h18a2, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hb553, 16'hb532, 16'hb512, 16'hb532, 16'hb532, 16'hb532, 16'had12, 16'had12, 16'hb512, 16'hb512, 16'hb532, 16'h944f, 16'h62a9, 16'h942e, 16'ha490, 16'h6ba, 16'h20e3, 16'h213, 16'h2923, 16'h18e2, 16'h840, 16'h840, 16'h840, 16'h860, 16'h841, 16'h840, 16'h860, 16'h840, 16'h840, 16'h840, 16'h840, 16'h840, 16'h841, 16'h1061, 16'h10a2, 16'h841, 16'h3964, 16'h6ac9, 16'h72e9, 16'h72e9, 16'h72e9, 16'h7ba, 16'h739, 16'h293, 16'h841, 16'h1882, 16'h293, 16'h293, 16'h62a8, 16'h6aa9, 16'h6aa9, 16'h72aa, 16'hb4d2, 16'hacb1, 16'h9cf, 16'hb4d2, 16'hb4d2, 16'hbd53, 16'h94f, 16'h8bad, 16'h4a7, 16'h3124, 16'h293, 16'h293, 16'h18a2, 16'h1081, 16'h18a2, 16'h214, 16'h841, 16'h820, 16'h292, 16'h41a3, 16'h41a4, 16'h41a4, 16'h3963, 16'h20e2, 16'h20e2, 16'h20e2, 16'h293, 16'h4a6, 16'h6aa9, 16'h73a, 16'h41a4, 16'h3984, 16'h3984, 16'h3964, 16'h3163, 16'h3163, 16'h3163, 16'h3164, 16'h213, 16'h840, 16'h820, 16'h820, 16'h820, 16'h820, 16'h820, 16'h840, 16'h20c1, 16'h3943, 16'h3943, 16'h3943, 16'h3943, 16'h3942, 16'h3943, 16'h3942, 16'h4184, 16'h3985, 16'h62aa, 16'hb532, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hb4d2, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d2, 16'hb4d1, 16'hb4f1, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb512, 16'hb4f2, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'h4a7, 16'h293, 16'h293, 16'h20e3, 16'h20e2, 16'h18a2, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hb553, 16'hbd53, 16'hb533, 16'hb533, 16'hb532, 16'hb532, 16'hb532, 16'hb512, 16'hb512, 16'had12, 16'hb512, 16'h942f, 16'h62a9, 16'h942f, 16'ha490, 16'h942e, 16'h838c, 16'h83ad, 16'h5267, 16'h20e2, 16'h860, 16'h860, 16'h860, 16'h860, 16'h860, 16'h860, 16'h860, 16'h860, 16'h840, 16'h840, 16'h861, 16'h2964, 16'h213, 16'h840, 16'h840, 16'h840, 16'h3964, 16'h6ac9, 16'h72e9, 16'h72e9, 16'h72ea, 16'h732a, 16'h739, 16'h293, 16'h841, 16'h841, 16'h18c5, 16'h20e5, 16'h6289, 16'h6aa9, 16'h6aa9, 16'h6269, 16'hb512, 16'hbd73, 16'h9c6f, 16'ha490, 16'hb4d2, 16'hbd33, 16'h94f, 16'h8bad, 16'h49e6, 16'h3164, 16'h3144, 16'h213, 16'h18a2, 16'h1081, 16'h18c2, 16'h2124, 16'h841, 16'h820, 16'h292, 16'h3984, 16'h41a4, 16'h41a4, 16'h41a4, 16'h3963, 16'h3123, 16'h2923, 16'h3143, 16'h5226, 16'h6aa8, 16'h73a, 16'h41c4, 16'h3984, 16'h3984, 16'h3963, 16'h3164, 16'h3164, 16'h3164, 16'h3984, 16'h3144, 16'h841, 16'h841, 16'h841, 16'h841, 16'h861, 16'h841, 16'h1061, 16'h20c1, 16'h3943, 16'h3943, 16'h3943, 16'h3943, 16'h3942, 16'h3943, 16'h3942, 16'h4164, 16'h3985, 16'h62ca, 16'hb512, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hacd2, 16'h4a7, 16'h293, 16'h212, 16'h20e2, 16'h20e2, 16'h18a1, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hb553, 16'hb532, 16'hb532, 16'hb532, 16'hb532, 16'hb532, 16'had12, 16'had12, 16'had12, 16'had12, 16'had12, 16'hb512, 16'h94e, 16'h62a9, 16'h942e, 16'ha4b0, 16'ha490, 16'h9c8f, 16'h9c4f, 16'h5a88, 16'h213, 16'h860, 16'h840, 16'h840, 16'h840, 16'h841, 16'h840, 16'h840, 16'h840, 16'h840, 16'h840, 16'h861, 16'h2944, 16'h20e3, 16'h840, 16'h840, 16'h820, 16'h3964, 16'h6ac9, 16'h72e9, 16'h72e9, 16'h72ea, 16'h7ba, 16'h72e9, 16'h293, 16'h841, 16'h296, 16'h3ad, 16'h31ab, 16'h62aa, 16'h6aa9, 16'h6aa9, 16'h6aca, 16'ha470, 16'hcdb5, 16'hb4f2, 16'h9c4f, 16'hacb1, 16'hbd33, 16'h93ee, 16'h838d, 16'h49e6, 16'h3164, 16'h3123, 16'h213, 16'h18c2, 16'h1081, 16'h18a2, 16'h213, 16'h841, 16'h820, 16'h292, 16'h3983, 16'h4184, 16'h3983, 16'h3963, 16'h3143, 16'h292, 16'h212, 16'h2923, 16'h49e5, 16'h6288, 16'h73a, 16'h41a4, 16'h3984, 16'h3984, 16'h3163, 16'h3163, 16'h3163, 16'h3163, 16'h3163, 16'h2923, 16'h840, 16'h020, 16'h820, 16'h820, 16'h840, 16'h840, 16'h1061, 16'h20e2, 16'h3143, 16'h3943, 16'h3943, 16'h3943, 16'h3942, 16'h3143, 16'h3142, 16'h3963, 16'h3985, 16'h62ca, 16'hb512, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f2, 16'hb4f2, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hacd2, 16'h4a7, 16'h293, 16'h212, 16'h20e2, 16'h20e2, 16'h18a1, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'hbd52, 16'hb552, 16'hbd53, 16'hbd53, 16'hb553, 16'hb552, 16'hb532, 16'hb532, 16'hb532, 16'had32, 16'had12, 16'had12, 16'had12, 16'had12, 16'had12, 16'had12, 16'h8ce, 16'h62a9, 16'h942e, 16'ha490, 16'ha490, 16'h9c6f, 16'h9c4e, 16'h5a88, 16'h212, 16'h860, 16'h840, 16'h840, 16'h840, 16'h860, 16'h860, 16'h840, 16'h840, 16'h840, 16'h840, 16'h840, 16'h840, 16'h840, 16'h840, 16'h840, 16'h841, 16'h3984, 16'h6ac9, 16'h72e9, 16'h72e9, 16'h72e9, 16'h7ba, 16'h6ae9, 16'h293, 16'h4a48, 16'h62ec, 16'h318b, 16'h3a2e, 16'h6bc, 16'h6aa9, 16'h62a9, 16'h7b2b, 16'h8bce, 16'hbd74, 16'hcdb5, 16'h94f, 16'ha491, 16'hb513, 16'h93ee, 16'h7b2b, 16'h3985, 16'h3965, 16'h3164, 16'h293, 16'h18c2, 16'h1061, 16'h18a2, 16'h213, 16'h841, 16'h820, 16'h292, 16'h41a4, 16'h41a4, 16'h4184, 16'h41a5, 16'h3964, 16'h2922, 16'h20e2, 16'h20e2, 16'h3143, 16'h41a5, 16'h5a47, 16'h41a4, 16'h3984, 16'h3984, 16'h3164, 16'h3163, 16'h3163, 16'h3164, 16'h2923, 16'h20e3, 16'h841, 16'h820, 16'h820, 16'h840, 16'h840, 16'h840, 16'h860, 16'h20e2, 16'h3143, 16'h3143, 16'h3143, 16'h3143, 16'h3143, 16'h3143, 16'h2923, 16'h3143, 16'h3164, 16'h5a89, 16'hb512, 16'hbd53, 16'hbd53, 16'hbd33, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hacf1, 16'hacf1, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hb4d1, 16'hb4d2, 16'hb4d2, 16'hb4d2, 16'hb4d2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb512, 16'hb4f2, 16'hacd2, 16'h4a7, 16'h293, 16'h20e2, 16'h20e2, 16'h20e2, 16'h18a1, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'hb532, 16'hb532, 16'hb552, 16'hb553, 16'hb553, 16'had32, 16'had12, 16'hb532, 16'had32, 16'had32, 16'hb532, 16'hb512, 16'had11, 16'had12, 16'had12, 16'had12, 16'h8bed, 16'h62a9, 16'h942e, 16'h94d, 16'h93ac, 16'h8b8b, 16'h8b6a, 16'h5227, 16'h212, 16'h840, 16'h840, 16'h840, 16'h840, 16'h860, 16'h840, 16'h841, 16'h840, 16'h840, 16'h840, 16'h020, 16'h020, 16'h020, 16'h840, 16'h861, 16'h861, 16'h3984, 16'h6ac9, 16'h6ac9, 16'h6ac9, 16'h6ac9, 16'h73a, 16'h6ac9, 16'h293, 16'h62eb, 16'h84f, 16'h2149, 16'h29ac, 16'h6aeb, 16'h6aa9, 16'h6aa9, 16'h7b2b, 16'h8bcd, 16'ha491, 16'hc5b5, 16'h93ee, 16'hacb1, 16'hb512, 16'h93ce, 16'h732b, 16'h3964, 16'h3144, 16'h3964, 16'h2923, 16'h18c2, 16'h1081, 16'h18a1, 16'h20e3, 16'h841, 16'h820, 16'h292, 16'h41a4, 16'h41a4, 16'h41c5, 16'h5247, 16'h4a6, 16'h39a4, 16'h3984, 16'h3984, 16'h49e6, 16'h5227, 16'h5a88, 16'h41a4, 16'h3984, 16'h3983, 16'h3163, 16'h3163, 16'h3163, 16'h3163, 16'h3143, 16'h213, 16'h18a2, 16'h10a2, 16'h10a1, 16'h10a1, 16'h18a1, 16'h10a2, 16'h10a1, 16'h18c2, 16'h20e2, 16'h18a1, 16'h18a1, 16'h1081, 16'h1081, 16'h1081, 16'h1081, 16'h1081, 16'h1881, 16'h4a7, 16'hb512, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hacf1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hb4d1, 16'hb4d2, 16'hb4d2, 16'hb4d2, 16'hb4d2, 16'hb4d2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hacb1, 16'h49e7, 16'h293, 16'h212, 16'h20e2, 16'h20e2, 16'h18a1, 16'h820, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'hb552, 16'hbd53, 16'hbd53, 16'hbd53, 16'hb533, 16'hb532, 16'had12, 16'hb532, 16'had32, 16'had12, 16'hb512, 16'hb512, 16'ha4f1, 16'ha4f2, 16'had12, 16'had12, 16'h83cd, 16'h62a9, 16'h942e, 16'h93cc, 16'h82e8, 16'h7ae7, 16'h7ac7, 16'h526, 16'h213, 16'h840, 16'h840, 16'h840, 16'h840, 16'h840, 16'h840, 16'h840, 16'h840, 16'h840, 16'h840, 16'h020, 16'h020, 16'h020, 16'h840, 16'h840, 16'h840, 16'h3144, 16'h5227, 16'h4a6, 16'h41c6, 16'h39a5, 16'h3984, 16'h3164, 16'h1081, 16'h2945, 16'h39c7, 16'h10a6, 16'h214b, 16'h62cb, 16'h6aa9, 16'h73b, 16'h836c, 16'h9cf, 16'h8bcf, 16'hacb2, 16'h93ce, 16'hb4f2, 16'hb4f2, 16'h8bad, 16'h732b, 16'h41a5, 16'h3144, 16'h3144, 16'h213, 16'h18c2, 16'h1081, 16'h18c2, 16'h18e2, 16'h840, 16'h020, 16'h18c2, 16'h2923, 16'h2944, 16'h2944, 16'h3965, 16'h49e6, 16'h49e6, 16'h49e6, 16'h4a7, 16'h5a48, 16'h72ea, 16'h73a, 16'h39a4, 16'h3984, 16'h3983, 16'h3163, 16'h3163, 16'h3163, 16'h3163, 16'h2923, 16'h20e2, 16'h1081, 16'h860, 16'h840, 16'h840, 16'h840, 16'h840, 16'h840, 16'h10a1, 16'h1081, 16'h860, 16'h860, 16'h860, 16'h860, 16'h860, 16'h860, 16'h1060, 16'h1081, 16'h41e6, 16'hb512, 16'hbd33, 16'hbd33, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd12, 16'hbd32, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f2, 16'hb4f1, 16'hacd1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hb4d2, 16'hb4d2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'ha4b1, 16'h4a7, 16'h293, 16'h212, 16'h20e2, 16'h20e2, 16'h18a2, 16'h820, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'had32, 16'hb532, 16'hbd52, 16'hbd52, 16'hb533, 16'hb532, 16'hb532, 16'hb532, 16'hb532, 16'hb532, 16'hb512, 16'had12, 16'ha4f1, 16'ha4f1, 16'hacf2, 16'had12, 16'h83cd, 16'h62a9, 16'h942e, 16'h9cc, 16'h624, 16'h4963, 16'h4983, 16'h41a5, 16'h213, 16'h860, 16'h840, 16'h840, 16'h861, 16'h860, 16'h860, 16'h860, 16'h860, 16'h860, 16'h860, 16'h840, 16'h840, 16'h840, 16'h840, 16'h840, 16'h840, 16'h861, 16'h861, 16'h861, 16'h840, 16'h840, 16'h840, 16'h840, 16'h040, 16'h020, 16'h040, 16'h042, 16'h18c5, 16'h62a9, 16'h6aa9, 16'h73b, 16'h73b, 16'h9c4f, 16'h9c30, 16'ha450, 16'ha470, 16'hb512, 16'hacb1, 16'h8bad, 16'h62a9, 16'h41c6, 16'h3985, 16'h3144, 16'h213, 16'h20e2, 16'h1081, 16'h18a2, 16'h18c2, 16'h841, 16'h020, 16'h1081, 16'h20e3, 16'h213, 16'h2924, 16'h3164, 16'h41a5, 16'h41a5, 16'h41c5, 16'h4a6, 16'h5247, 16'h6ac9, 16'h6ae9, 16'h39a4, 16'h3984, 16'h3163, 16'h3163, 16'h3164, 16'h3163, 16'h3164, 16'h2923, 16'h20e2, 16'h1081, 16'h840, 16'h840, 16'h840, 16'h840, 16'h840, 16'h860, 16'h18a1, 16'h1061, 16'h860, 16'h860, 16'h1060, 16'h1080, 16'h1081, 16'h1081, 16'h1081, 16'h18a1, 16'h4a6, 16'hb512, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f2, 16'hb4f2, 16'hacf2, 16'hacf1, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacd1, 16'hacb1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hb4d2, 16'hb4d1, 16'hb4d2, 16'hb4d2, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hb4f1, 16'hb4f2, 16'hb4f2, 16'ha490, 16'h49e6, 16'h213, 16'h212, 16'h20e2, 16'h20e2, 16'h18a1, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'hb532, 16'hb532, 16'hb532, 16'hb532, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'had12, 16'had12, 16'ha4f1, 16'ha4f1, 16'hacf2, 16'had12, 16'h83ad, 16'h62a9, 16'h942e, 16'h9bec, 16'h4983, 16'h3922, 16'h3942, 16'h39c5, 16'h2123, 16'h840, 16'h840, 16'h861, 16'h18c2, 16'h861, 16'h860, 16'h840, 16'h840, 16'h840, 16'h040, 16'h040, 16'h040, 16'h040, 16'h840, 16'h840, 16'h840, 16'h040, 16'h040, 16'h040, 16'h840, 16'h840, 16'h040, 16'h840, 16'h040, 16'h020, 16'h840, 16'h841, 16'h1082, 16'h62a8, 16'h6ac9, 16'h6289, 16'h4186, 16'h8bad, 16'hb4f2, 16'hb4f2, 16'hb512, 16'hb4f2, 16'ha470, 16'h8b8d, 16'h5a48, 16'h3985, 16'h39a5, 16'h3964, 16'h2924, 16'h213, 16'h1081, 16'h18a2, 16'h18c2, 16'h840, 16'h020, 16'h1081, 16'h20c2, 16'h3144, 16'h41a5, 16'h41c5, 16'h41c5, 16'h41a5, 16'h49e6, 16'h49e6, 16'h41a5, 16'h526, 16'h62a8, 16'h39a4, 16'h3984, 16'h3163, 16'h3163, 16'h3163, 16'h3164, 16'h3164, 16'h3143, 16'h213, 16'h1061, 16'h860, 16'h860, 16'h861, 16'h1081, 16'h1081, 16'h18a2, 16'h18c1, 16'h1081, 16'h10a1, 16'h10a1, 16'h18c1, 16'h18c1, 16'h18c1, 16'h18c2, 16'h18e2, 16'h212, 16'h5247, 16'hb512, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f2, 16'hacf1, 16'hacf1, 16'hacf1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hb4d1, 16'hb4d1, 16'ha490, 16'h4a6, 16'h293, 16'h212, 16'h20e2, 16'h20e2, 16'h18a1, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'hb532, 16'hb532, 16'had12, 16'hb532, 16'hb4f2, 16'hacf2, 16'hacf2, 16'hacf1, 16'hb512, 16'hb512, 16'had12, 16'hacf2, 16'ha4d1, 16'hacf1, 16'hacf2, 16'hacf1, 16'h838c, 16'h62a9, 16'h942e, 16'h9bec, 16'h51a3, 16'h392, 16'h3122, 16'h39a5, 16'h2123, 16'h840, 16'h840, 16'h861, 16'h18e3, 16'h861, 16'h840, 16'h840, 16'h840, 16'h840, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h020, 16'h040, 16'h840, 16'h840, 16'h1081, 16'h6288, 16'h6ac9, 16'h6ac9, 16'h527, 16'h73b, 16'hb4f2, 16'hb4f2, 16'hacd1, 16'hb4f2, 16'h9cf, 16'h838d, 16'h4a6, 16'h3964, 16'h41a5, 16'h41a6, 16'h2944, 16'h2123, 16'h1081, 16'h18a2, 16'h18a2, 16'h840, 16'h020, 16'h1081, 16'h20e2, 16'h3164, 16'h41a5, 16'h41a5, 16'h41c5, 16'h41a4, 16'h4a6, 16'h6ac8, 16'h5a67, 16'h526, 16'h5a67, 16'h39a4, 16'h3983, 16'h3183, 16'h3163, 16'h3963, 16'h3164, 16'h3164, 16'h3164, 16'h2923, 16'h18a1, 16'h10a1, 16'h18c1, 16'h18c2, 16'h18c2, 16'h18e2, 16'h18e2, 16'h18e2, 16'h20e2, 16'h20e2, 16'h212, 16'h212, 16'h212, 16'h213, 16'h2123, 16'h2923, 16'h2943, 16'h5268, 16'hb4f2, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hbd32, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hacd1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'h9c6f, 16'h41c6, 16'h293, 16'h212, 16'h20e2, 16'h20e2, 16'h18a1, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'hbd32, 16'hb532, 16'had12, 16'hb532, 16'hb512, 16'hb512, 16'hacf1, 16'hacf2, 16'hb512, 16'hb512, 16'had12, 16'hacf2, 16'ha4f1, 16'hacf1, 16'hacf1, 16'hacf1, 16'h838c, 16'h62a9, 16'h94e, 16'h9beb, 16'h4983, 16'h311, 16'h3122, 16'h41c5, 16'h2944, 16'h840, 16'h840, 16'h861, 16'h213, 16'h10a2, 16'h040, 16'h840, 16'h840, 16'h840, 16'h040, 16'h040, 16'h840, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h020, 16'h020, 16'h020, 16'h040, 16'h840, 16'h840, 16'h1081, 16'h6288, 16'h6ac9, 16'h6ac9, 16'h6ac9, 16'h49e6, 16'h6aaa, 16'ha470, 16'hacb1, 16'hb512, 16'h8bcd, 16'h7b6c, 16'h41a5, 16'h3964, 16'h41c6, 16'h49e6, 16'h3144, 16'h2923, 16'h1081, 16'h18a2, 16'h18a2, 16'h840, 16'h020, 16'h861, 16'h1881, 16'h20e2, 16'h3143, 16'h3143, 16'h3143, 16'h2923, 16'h2943, 16'h41a4, 16'h4a5, 16'h49e6, 16'h5226, 16'h3984, 16'h3984, 16'h3983, 16'h3963, 16'h3963, 16'h3963, 16'h3163, 16'h3143, 16'h20e2, 16'h20e2, 16'h212, 16'h212, 16'h212, 16'h212, 16'h213, 16'h213, 16'h2123, 16'h2123, 16'h2923, 16'h2923, 16'h2923, 16'h2943, 16'h2943, 16'h2943, 16'h2943, 16'h3164, 16'h5a68, 16'hb4f2, 16'hbd32, 16'hbd32, 16'hbd32, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hacd1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'h9c70, 16'h41c6, 16'h213, 16'h212, 16'h20e2, 16'h20e2, 16'h18a1, 16'h820, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'hbd52, 16'hb532, 16'hb532, 16'hb532, 16'hb532, 16'hb532, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hacf2, 16'hacf2, 16'ha4d1, 16'hacf1, 16'hacf1, 16'hacf1, 16'h7b6c, 16'h62a9, 16'h94e, 16'h9beb, 16'h4983, 16'h3121, 16'h3922, 16'h41c6, 16'h2944, 16'h840, 16'h860, 16'h861, 16'h213, 16'h18c2, 16'h841, 16'h040, 16'h840, 16'h040, 16'h040, 16'h840, 16'h840, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h840, 16'h840, 16'h1081, 16'h6287, 16'h6ac9, 16'h6ac9, 16'h6ac9, 16'h6288, 16'h4185, 16'h6289, 16'h9c70, 16'hacb1, 16'h838d, 16'h73b, 16'h3964, 16'h3985, 16'h5227, 16'h5227, 16'h3144, 16'h2944, 16'h20e2, 16'h20e2, 16'h18c2, 16'h840, 16'h020, 16'h1061, 16'h20c2, 16'h212, 16'h292, 16'h292, 16'h292, 16'h292, 16'h2923, 16'h2943, 16'h2923, 16'h20e2, 16'h39a4, 16'h3984, 16'h3984, 16'h3983, 16'h3984, 16'h3964, 16'h3163, 16'h3163, 16'h3143, 16'h2123, 16'h2123, 16'h2123, 16'h2123, 16'h2123, 16'h2923, 16'h2923, 16'h2923, 16'h2923, 16'h2923, 16'h2923, 16'h2923, 16'h2943, 16'h2943, 16'h2943, 16'h2944, 16'h3144, 16'h3164, 16'h5a68, 16'hb4f1, 16'hbd32, 16'hbd32, 16'hbd32, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacd1, 16'hacb1, 16'h9c2f, 16'h49e6, 16'h293, 16'h212, 16'h20e2, 16'h20e2, 16'h18c1, 16'h820, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'hbd52, 16'hbd32, 16'hb532, 16'hb532, 16'hb532, 16'hb532, 16'hb512, 16'hb512, 16'hb512, 16'hacf2, 16'hacd1, 16'hacd1, 16'ha4d1, 16'hacd1, 16'ha4d1, 16'hacd1, 16'h7b6b, 16'h62a9, 16'h94e, 16'h93ca, 16'h4962, 16'h30e1, 16'h3922, 16'h526, 16'h3144, 16'h840, 16'h860, 16'h861, 16'h213, 16'h18e2, 16'h861, 16'h020, 16'h040, 16'h040, 16'h040, 16'h840, 16'h840, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h840, 16'h840, 16'h840, 16'h840, 16'h1081, 16'h6288, 16'h6ac9, 16'h6ac9, 16'h6ac9, 16'h6ac9, 16'h6288, 16'h49c6, 16'h62aa, 16'h8bce, 16'h7b2b, 16'h5a68, 16'h3144, 16'h41a5, 16'h5a48, 16'h5a68, 16'h3144, 16'h39a5, 16'h4a6, 16'h213, 16'h18c2, 16'h841, 16'h020, 16'h1061, 16'h18c2, 16'h18c1, 16'h20c2, 16'h20e2, 16'h20e2, 16'h20e2, 16'h20c1, 16'h20c1, 16'h18c2, 16'h212, 16'h3984, 16'h3984, 16'h3984, 16'h3984, 16'h3984, 16'h3143, 16'h3143, 16'h3143, 16'h2923, 16'h212, 16'h2123, 16'h2123, 16'h2923, 16'h2123, 16'h2923, 16'h2923, 16'h2943, 16'h2923, 16'h2923, 16'h2943, 16'h2943, 16'h2943, 16'h2943, 16'h2943, 16'h2944, 16'h3164, 16'h3164, 16'h5a68, 16'hb4f2, 16'hbd32, 16'hbd32, 16'hbd32, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'ha490, 16'hacb0, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'ha4b0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'h9c4f, 16'h49e7, 16'h293, 16'h212, 16'h20e2, 16'h20e2, 16'h18a1, 16'h820, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'hb532, 16'hb532, 16'hb532, 16'hb532, 16'hb532, 16'hb512, 16'hb512, 16'hb512, 16'hacf2, 16'hacf1, 16'ha4d0, 16'ha4d1, 16'ha4d1, 16'ha4d1, 16'ha4b1, 16'hacd0, 16'h7b4b, 16'h62a9, 16'h94e, 16'h93aa, 16'h4162, 16'h30e1, 16'h3122, 16'h4a6, 16'h3164, 16'h840, 16'h040, 16'h861, 16'h18e2, 16'h18c2, 16'h1061, 16'h020, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h841, 16'h861, 16'h1061, 16'h840, 16'h1081, 16'h6267, 16'h6ac9, 16'h6ac9, 16'h6ac9, 16'h6ac9, 16'h6ac9, 16'h6aa9, 16'h6aca, 16'h5a89, 16'h3144, 16'h20e3, 16'h18a2, 16'h3144, 16'h4a7, 16'h5227, 16'h41a6, 16'h4a7, 16'h5248, 16'h20e2, 16'h18c2, 16'h841, 16'h020, 16'h1061, 16'h18c2, 16'h20e2, 16'h20e3, 16'h293, 16'h213, 16'h213, 16'h213, 16'h212, 16'h20e2, 16'h20e2, 16'h3984, 16'h39a4, 16'h39a4, 16'h3984, 16'h3963, 16'h2922, 16'h2923, 16'h2943, 16'h2923, 16'h2123, 16'h2123, 16'h2123, 16'h2123, 16'h2923, 16'h2923, 16'h2923, 16'h2923, 16'h2943, 16'h2923, 16'h2943, 16'h2943, 16'h2943, 16'h2943, 16'h2943, 16'h2944, 16'h3143, 16'h3144, 16'h5a68, 16'hb4f1, 16'hbd32, 16'hbd32, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'ha490, 16'ha490, 16'hacb0, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'ha4b0, 16'ha4b0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'ha4b0, 16'hacb0, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'ha4b0, 16'ha4b0, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'h9c2f, 16'h49e6, 16'h293, 16'h212, 16'h20e2, 16'h20e2, 16'h18c1, 16'h820, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'hb532, 16'hb512, 16'hb532, 16'hb532, 16'hb532, 16'hb512, 16'hb512, 16'hb512, 16'hacf2, 16'hacf1, 16'ha4d1, 16'ha4d0, 16'ha4b0, 16'ha4b0, 16'ha4b0, 16'ha4d0, 16'h734b, 16'h62a9, 16'h94d, 16'h93aa, 16'h4962, 16'h312, 16'h3122, 16'h4a6, 16'h2944, 16'h840, 16'h040, 16'h861, 16'h20e2, 16'h18c2, 16'h1081, 16'h020, 16'h020, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h020, 16'h020, 16'h020, 16'h020, 16'h860, 16'h861, 16'h840, 16'h10a2, 16'h1881, 16'h840, 16'h1081, 16'h6267, 16'h6ac9, 16'h6ac9, 16'h6ac9, 16'h6ac9, 16'h6ae9, 16'h72e9, 16'h7b2b, 16'h3985, 16'h1881, 16'h18c2, 16'h18a2, 16'h20e3, 16'h2923, 16'h293, 16'h3985, 16'h4a27, 16'h5227, 16'h20c2, 16'h1081, 16'h840, 16'h020, 16'h1081, 16'h213, 16'h213, 16'h213, 16'h213, 16'h213, 16'h213, 16'h3184, 16'h41c5, 16'h41a5, 16'h2923, 16'h3964, 16'h39a4, 16'h3984, 16'h3964, 16'h3163, 16'h3143, 16'h3143, 16'h3143, 16'h2923, 16'h213, 16'h213, 16'h213, 16'h213, 16'h212, 16'h213, 16'h213, 16'h213, 16'h2923, 16'h2923, 16'h2943, 16'h2943, 16'h3143, 16'h3164, 16'h3164, 16'h3184, 16'h3984, 16'h3984, 16'h5a88, 16'hb4f1, 16'hb532, 16'hbd32, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'ha490, 16'ha490, 16'hac90, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'ha4b0, 16'ha4b0, 16'ha490, 16'hac90, 16'hac90, 16'hacb0, 16'hacb0, 16'hacb0, 16'ha4b0, 16'ha4b0, 16'ha4b0, 16'ha4b0, 16'hacb1, 16'hacb0, 16'ha4b0, 16'ha490, 16'ha4b0, 16'hacb0, 16'hacb0, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'ha4b1, 16'ha490, 16'h9c2f, 16'h49e6, 16'h293, 16'h212, 16'h20e2, 16'h20e2, 16'h18c1, 16'h820, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'hb511, 16'hb512, 16'hb512, 16'hb512, 16'hb532, 16'hb512, 16'hb512, 16'hb512, 16'hacf1, 16'hacf1, 16'hacf1, 16'ha4d1, 16'ha4d1, 16'ha4d1, 16'ha4d0, 16'ha4b0, 16'h732b, 16'h62a9, 16'h7b6b, 16'h8b89, 16'h4162, 16'h30e1, 16'h312, 16'h4a26, 16'h213, 16'h040, 16'h040, 16'h861, 16'h20e3, 16'h18e2, 16'h1081, 16'h020, 16'h020, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h820, 16'h840, 16'h18c2, 16'h18a2, 16'h840, 16'h1061, 16'h6267, 16'h6ac9, 16'h6ac9, 16'h6ac9, 16'h6ac9, 16'h6ae9, 16'h72e9, 16'h6ac9, 16'h41c5, 16'h20e2, 16'h820, 16'h840, 16'h820, 16'h820, 16'h020, 16'h841, 16'h18a2, 16'h3144, 16'h20e3, 16'h1081, 16'h840, 16'h020, 16'h2944, 16'h5227, 16'h3184, 16'h31a4, 16'h18c2, 16'h1061, 16'h18a2, 16'h62a8, 16'h7b6b, 16'h732a, 16'h4a6, 16'h41a5, 16'h39a4, 16'h3984, 16'h3163, 16'h3143, 16'h3142, 16'h2943, 16'h2943, 16'h2923, 16'h2122, 16'h2923, 16'h2923, 16'h2943, 16'h3163, 16'h3163, 16'h3164, 16'h3164, 16'h3164, 16'h3184, 16'h3164, 16'h3164, 16'h3164, 16'h3984, 16'h3964, 16'h3984, 16'h3964, 16'h3984, 16'h5a68, 16'hb4f1, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'ha4b0, 16'hacb0, 16'ha4b0, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'hac90, 16'ha490, 16'ha490, 16'hacb0, 16'ha4b0, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha4b0, 16'ha4b0, 16'ha4b0, 16'ha490, 16'ha4b0, 16'ha4b0, 16'ha4b0, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha4b0, 16'ha4b0, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'ha490, 16'ha490, 16'h942e, 16'h49e6, 16'h293, 16'h212, 16'h20e2, 16'h20e2, 16'h18c1, 16'h820, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'hacf1, 16'hacf1, 16'hb4f1, 16'hb511, 16'hb511, 16'hb512, 16'hb512, 16'hb512, 16'hacf1, 16'hacf1, 16'hacf1, 16'ha4d1, 16'ha4b0, 16'ha4b0, 16'ha490, 16'h9c6f, 16'h732a, 16'h62a9, 16'h5a47, 16'h7ac7, 16'h4122, 16'h28c1, 16'h30e2, 16'h49e6, 16'h18c2, 16'h840, 16'h840, 16'h1081, 16'h213, 16'h18e2, 16'h881, 16'h020, 16'h020, 16'h020, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h840, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h820, 16'h840, 16'h861, 16'h840, 16'h820, 16'h1081, 16'h6287, 16'h6ac9, 16'h6ac9, 16'h6ac9, 16'h6ac9, 16'h6ae9, 16'h72e9, 16'h7b2a, 16'h6ac8, 16'h2923, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h841, 16'h1061, 16'h1061, 16'h820, 16'h820, 16'h5268, 16'h9c6f, 16'h4a47, 16'h52c8, 16'h2964, 16'h861, 16'h1061, 16'h39a5, 16'h39a5, 16'h2924, 16'h20e3, 16'h41a4, 16'h3163, 16'h3163, 16'h3143, 16'h2942, 16'h2922, 16'h212, 16'h2922, 16'h2942, 16'h2943, 16'h2943, 16'h2943, 16'h3143, 16'h3143, 16'h3143, 16'h3143, 16'h3143, 16'h3143, 16'h3143, 16'h3143, 16'h3143, 16'h3143, 16'h3164, 16'h3163, 16'h3163, 16'h3163, 16'h3964, 16'h5a68, 16'hb4f1, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'ha4b0, 16'ha490, 16'ha490, 16'ha490, 16'hac90, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha4b0, 16'ha4b0, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha4b0, 16'ha4b0, 16'ha4b0, 16'ha4b1, 16'hacb1, 16'ha4b1, 16'ha4b0, 16'ha491, 16'ha491, 16'ha490, 16'h94e, 16'h49e6, 16'h293, 16'h212, 16'h212, 16'h20e2, 16'h18c1, 16'h820, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'ha4af, 16'ha4b0, 16'ha4b0, 16'ha4b0, 16'ha4b0, 16'ha4b0, 16'ha4b0, 16'ha490, 16'h9c70, 16'h9c6f, 16'h9c4f, 16'h944f, 16'h942e, 16'h942e, 16'h94e, 16'h94e, 16'h83cd, 16'h83ac, 16'h6288, 16'h7ae8, 16'h3921, 16'h30e1, 16'h391, 16'h4163, 16'h3122, 16'h3121, 16'h3942, 16'h4183, 16'h3163, 16'h20e2, 16'h1081, 16'h020, 16'h020, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h840, 16'h840, 16'h840, 16'h020, 16'h020, 16'h020, 16'h020, 16'h861, 16'h2123, 16'h1081, 16'h020, 16'h020, 16'h020, 16'h020, 16'h1081, 16'h6288, 16'h6ac9, 16'h6ac9, 16'h6ac9, 16'h6ac9, 16'h6ac9, 16'h72e9, 16'h7b4a, 16'h6ac9, 16'h293, 16'h820, 16'h820, 16'h840, 16'h841, 16'h840, 16'h840, 16'h840, 16'h840, 16'h840, 16'h861, 16'h840, 16'h020, 16'h49e7, 16'ha490, 16'h39a6, 16'h39e5, 16'h3184, 16'h861, 16'h840, 16'h820, 16'h020, 16'h020, 16'h840, 16'h20c2, 16'h18c1, 16'h20e1, 16'h211, 16'h20e2, 16'h18c1, 16'h18c1, 16'h212, 16'h212, 16'h2122, 16'h2922, 16'h2922, 16'h2922, 16'h2922, 16'h2923, 16'h2923, 16'h2923, 16'h2923, 16'h2922, 16'h292, 16'h212, 16'h20e2, 16'h20e2, 16'h20e2, 16'h20e2, 16'h20c2, 16'h20c2, 16'h49e7, 16'hacd1, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'ha4b0, 16'ha4b0, 16'ha490, 16'hac90, 16'ha490, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha4b0, 16'ha4b0, 16'ha4b0, 16'ha4b0, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha4b0, 16'ha4b0, 16'hac91, 16'hac91, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'h94e, 16'h49e6, 16'h293, 16'h212, 16'h20e2, 16'h20e2, 16'h18c1, 16'h820, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h8bcd, 16'h93ed, 16'h94e, 16'h942e, 16'h9c4e, 16'h9c4f, 16'h9c6f, 16'h9c6f, 16'h9c70, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'h9c90, 16'h9c6f, 16'h9c4f, 16'h942e, 16'h6288, 16'h7ac7, 16'h4962, 16'h4141, 16'h4962, 16'h51a3, 16'h59c3, 16'h59e3, 16'h59e4, 16'h6a66, 16'h3984, 16'h20c2, 16'h1081, 16'h020, 16'h040, 16'h020, 16'h040, 16'h020, 16'h840, 16'h840, 16'h840, 16'h840, 16'h840, 16'h020, 16'h020, 16'h020, 16'h020, 16'h18c2, 16'h4a47, 16'h18c2, 16'h020, 16'h020, 16'h820, 16'h841, 16'h1882, 16'h6288, 16'h6ac9, 16'h6ac9, 16'h6ac9, 16'h6ac9, 16'h6ac9, 16'h72e9, 16'h7b4a, 16'h6ac8, 16'h3144, 16'h18c2, 16'h18c2, 16'h18c2, 16'h10a2, 16'h1081, 16'h10a2, 16'h10a2, 16'h1081, 16'h1081, 16'h18a2, 16'h10a2, 16'h020, 16'h20e3, 16'h6aea, 16'h2924, 16'h861, 16'h840, 16'h020, 16'h020, 16'h841, 16'h861, 16'h841, 16'h1061, 16'h20e2, 16'h20e1, 16'h20e2, 16'h20e1, 16'h20e2, 16'h18c1, 16'h18c1, 16'h18c1, 16'h18c1, 16'h18c1, 16'h18a1, 16'h10a1, 16'h1081, 16'h1081, 16'h1081, 16'h1061, 16'h861, 16'h840, 16'h840, 16'h840, 16'h840, 16'h840, 16'h840, 16'h840, 16'h841, 16'h861, 16'h1061, 16'h41a6, 16'hacd1, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4d2, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'hac90, 16'hac90, 16'hac90, 16'ha4b0, 16'ha4b0, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha4b0, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'h94e, 16'h49e6, 16'h293, 16'h212, 16'h20e2, 16'h20e2, 16'h18c1, 16'h820, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h94d, 16'h942e, 16'h9c4f, 16'h9c6f, 16'ha490, 16'ha490, 16'ha490, 16'ha4b0, 16'ha4b0, 16'ha4b0, 16'ha4b0, 16'ha4b0, 16'ha490, 16'ha490, 16'ha490, 16'h9c6f, 16'h9c6f, 16'h942e, 16'h5247, 16'h525, 16'h4983, 16'h4163, 16'h3942, 16'h3922, 16'h312, 16'h28c2, 16'h3944, 16'h6ae9, 16'h41c5, 16'h20c2, 16'h1081, 16'h020, 16'h020, 16'h020, 16'h020, 16'h040, 16'h840, 16'h840, 16'h020, 16'h840, 16'h840, 16'h020, 16'h020, 16'h020, 16'h020, 16'h1081, 16'h3164, 16'h10a2, 16'h020, 16'h020, 16'h020, 16'h020, 16'h1081, 16'h6287, 16'h6ac9, 16'h6ac9, 16'h6ac9, 16'h6ac9, 16'h72e9, 16'h72e9, 16'h73a, 16'h5247, 16'h3164, 16'h2924, 16'h213, 16'h213, 16'h18c2, 16'h18c2, 16'h18c2, 16'h18a2, 16'h10a2, 16'h10a1, 16'h18a2, 16'h1081, 16'h020, 16'h020, 16'h1061, 16'h820, 16'h020, 16'h840, 16'h841, 16'h862, 16'h1083, 16'h1082, 16'h861, 16'h18a2, 16'h4185, 16'h5247, 16'h5a88, 16'h3143, 16'h18a1, 16'h841, 16'h840, 16'h840, 16'h840, 16'h840, 16'h820, 16'h840, 16'h840, 16'h840, 16'h840, 16'h840, 16'h860, 16'h861, 16'h1061, 16'h1081, 16'h1081, 16'h1081, 16'h10a1, 16'h10a1, 16'h10a1, 16'h1082, 16'h1882, 16'h41c6, 16'hacd1, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'ha490, 16'hac90, 16'hacb0, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha490, 16'ha470, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'h94e, 16'h49e6, 16'h213, 16'h212, 16'h20e2, 16'h20e2, 16'h18c1, 16'h820, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h8bcd, 16'h94d, 16'h942e, 16'h9c2f, 16'h9c4f, 16'h9c6f, 16'h9c70, 16'ha46f, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'h9c90, 16'h9c6f, 16'h9c6f, 16'h942e, 16'h4a26, 16'h18a2, 16'h860, 16'h860, 16'h840, 16'h840, 16'h840, 16'h840, 16'h3164, 16'h7b4b, 16'h41c6, 16'h20e2, 16'h1081, 16'h020, 16'h020, 16'h020, 16'h020, 16'h040, 16'h040, 16'h840, 16'h020, 16'h040, 16'h040, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h840, 16'h840, 16'h840, 16'h1081, 16'h6288, 16'h72c9, 16'h6ac9, 16'h72c9, 16'h72c9, 16'h72c9, 16'h6ac9, 16'h5248, 16'h3985, 16'h3144, 16'h2923, 16'h213, 16'h213, 16'h20e3, 16'h20e3, 16'h20e3, 16'h18e2, 16'h18c2, 16'h18c2, 16'h18c2, 16'h10a2, 16'h841, 16'h840, 16'h861, 16'h840, 16'h1881, 16'h18c2, 16'h18c3, 16'h20e4, 16'h215, 16'h2923, 16'h2923, 16'h3144, 16'h5227, 16'h72e9, 16'h8bcc, 16'h73a, 16'h39a4, 16'h20e2, 16'h861, 16'h840, 16'h840, 16'h040, 16'h020, 16'h840, 16'h840, 16'h840, 16'h840, 16'h840, 16'h861, 16'h1061, 16'h1061, 16'h1061, 16'h861, 16'h841, 16'h840, 16'h840, 16'h840, 16'h841, 16'h1061, 16'h4185, 16'hacd1, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'h9c50, 16'h93ee, 16'h49e6, 16'h212, 16'h212, 16'h212, 16'h20e2, 16'h18c1, 16'h820, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h838c, 16'h8bcc, 16'h8bed, 16'h94e, 16'h942e, 16'h942e, 16'h9c4f, 16'h9c4f, 16'h9c6f, 16'h9c6f, 16'h9c6f, 16'h9c70, 16'h9c70, 16'h9c6f, 16'h9c6f, 16'h9c6f, 16'h9c4f, 16'h942e, 16'h4a6, 16'h1081, 16'h840, 16'h040, 16'h040, 16'h040, 16'h840, 16'h840, 16'h2944, 16'h732b, 16'h41e6, 16'h18e2, 16'h1081, 16'h020, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h00, 16'h020, 16'h020, 16'h841, 16'h861, 16'h861, 16'h18a2, 16'h6288, 16'h6ac9, 16'h72c9, 16'h72c9, 16'h72c9, 16'h6ac9, 16'h5a68, 16'h39a6, 16'h3144, 16'h2924, 16'h2123, 16'h213, 16'h20e3, 16'h2124, 16'h2124, 16'h18e3, 16'h18c2, 16'h18c2, 16'h18e2, 16'h20e3, 16'h215, 16'h18a5, 16'h20c2, 16'h28e2, 16'h292, 16'h4184, 16'h49c5, 16'h41e6, 16'h4a6, 16'h527, 16'h4a6, 16'h4a6, 16'h4a6, 16'h5227, 16'h6288, 16'h838b, 16'ha48f, 16'h8bcd, 16'h5226, 16'h2923, 16'h861, 16'h020, 16'h020, 16'h020, 16'h020, 16'h820, 16'h820, 16'h820, 16'h840, 16'h840, 16'h840, 16'h840, 16'h840, 16'h840, 16'h840, 16'h1061, 16'h1061, 16'h1081, 16'h18a1, 16'h20c2, 16'h49e6, 16'hacd1, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hacb0, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha46f, 16'ha46f, 16'ha470, 16'ha470, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'h9c50, 16'h9c50, 16'h93ee, 16'h49e6, 16'h213, 16'h212, 16'h20e2, 16'h20e2, 16'h18c1, 16'h820, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h7b4b, 16'h7b6c, 16'h83ad, 16'h8bcd, 16'h8bed, 16'h94e, 16'h94e, 16'h942e, 16'h9c2f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h94e, 16'h426, 16'h1081, 16'h840, 16'h840, 16'h040, 16'h040, 16'h040, 16'h040, 16'h2944, 16'h734b, 16'h4a7, 16'h18c2, 16'h861, 16'h020, 16'h020, 16'h020, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h00, 16'h020, 16'h020, 16'h841, 16'h1081, 16'h861, 16'h1882, 16'h6288, 16'h72c9, 16'h72c9, 16'h72c9, 16'h72c9, 16'h6ac9, 16'h49e7, 16'h3165, 16'h2924, 16'h294, 16'h213, 16'h213, 16'h20e3, 16'h20e3, 16'h20e3, 16'h18e3, 16'h18e2, 16'h20e2, 16'h213, 16'h3165, 16'h2947, 16'h2128, 16'h28e3, 16'h3123, 16'h5247, 16'h5227, 16'h5227, 16'h5227, 16'h5227, 16'h5227, 16'h5227, 16'h4a6, 16'h49e5, 16'h49e6, 16'h5227, 16'h6aa9, 16'h8b8c, 16'hac90, 16'h93ed, 16'h5226, 16'h2943, 16'h840, 16'h820, 16'h840, 16'h841, 16'h861, 16'h1081, 16'h18a1, 16'h18a2, 16'h20c2, 16'h212, 16'h2923, 16'h3144, 16'h3164, 16'h3984, 16'h39a4, 16'h41c5, 16'h41e5, 16'h49e5, 16'h4a6, 16'h6aa9, 16'hacd1, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha46f, 16'ha46f, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha490, 16'ha490, 16'ha470, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'h9c6f, 16'h9c4f, 16'h9c4f, 16'h93ee, 16'h4a6, 16'h213, 16'h212, 16'h20e2, 16'h20e2, 16'h18c1, 16'h820, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h732a, 16'h7b2b, 16'h7b6b, 16'h838c, 16'h83ac, 16'h8bad, 16'h8bcd, 16'h93ee, 16'h94e, 16'h942e, 16'h942f, 16'h942f, 16'h942f, 16'h9c2e, 16'h9c2f, 16'h9c2f, 16'h942f, 16'h94e, 16'h41e5, 16'h1081, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h39a5, 16'h6bb, 16'h427, 16'h18e2, 16'h881, 16'h020, 16'h040, 16'h020, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h00, 16'h020, 16'h020, 16'h840, 16'h841, 16'h840, 16'h1881, 16'h6288, 16'h6ac9, 16'h6ac9, 16'h72c9, 16'h72c9, 16'h6288, 16'h41a5, 16'h3164, 16'h2923, 16'h213, 16'h20e3, 16'h213, 16'h20e3, 16'h20e3, 16'h20e2, 16'h20e2, 16'h20e2, 16'h20e3, 16'h41e7, 16'h7b8d, 16'h3986, 16'h2129, 16'h18c6, 16'h28e4, 16'h7b6c, 16'h838c, 16'h5227, 16'h5227, 16'h4a6, 16'h49e6, 16'h49e5, 16'h49c5, 16'h49c5, 16'h49e5, 16'h525, 16'h5a46, 16'h6a87, 16'h834a, 16'ha44e, 16'h6ac9, 16'h41e5, 16'h18c2, 16'h18c2, 16'h2922, 16'h3164, 16'h39a4, 16'h41c5, 16'h49e5, 16'h49e5, 16'h49e5, 16'h49e5, 16'h49e5, 16'h41c5, 16'h41c5, 16'h41a5, 16'h3984, 16'h3964, 16'h3164, 16'h3143, 16'h2923, 16'h527, 16'hacb1, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha44f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha46f, 16'ha470, 16'ha470, 16'ha470, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h93ee, 16'h4a6, 16'h213, 16'h212, 16'h20e2, 16'h20e2, 16'h18c1, 16'h820, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h6aea, 16'h73a, 16'h732a, 16'h7b4b, 16'h7b4b, 16'h838c, 16'h83ac, 16'h8bad, 16'h8bcd, 16'h8bed, 16'h93ed, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h942e, 16'h94e, 16'h8bed, 16'h41c5, 16'h881, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h10a2, 16'h31a6, 16'h4a27, 16'h18c2, 16'h1081, 16'h020, 16'h040, 16'h020, 16'h020, 16'h840, 16'h040, 16'h040, 16'h040, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h1061, 16'h6267, 16'h72c9, 16'h6ac9, 16'h6ac9, 16'h6ac9, 16'h5a47, 16'h3985, 16'h3144, 16'h2923, 16'h213, 16'h213, 16'h213, 16'h20e3, 16'h18c2, 16'h20e3, 16'h20e2, 16'h20e2, 16'h20e3, 16'h3986, 16'h942f, 16'h5a89, 16'h2949, 16'h214b, 16'h10a8, 16'h4a2b, 16'ha491, 16'h739, 16'h41a4, 16'h41a4, 16'h41a4, 16'h49c4, 16'h49c4, 16'h51e5, 16'h525, 16'h5a26, 16'h5a26, 16'h6267, 16'h72c8, 16'h93ed, 16'h6ac9, 16'h41e5, 16'h20e2, 16'h20e2, 16'h2923, 16'h3143, 16'h3143, 16'h2923, 16'h293, 16'h20e3, 16'h20c2, 16'h18a2, 16'h1881, 16'h1081, 16'h1061, 16'h861, 16'h840, 16'h840, 16'h840, 16'h840, 16'h840, 16'h3965, 16'hacb1, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hacb0, 16'hacb0, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha46f, 16'ha470, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha450, 16'ha46f, 16'ha46f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'ha46f, 16'ha470, 16'ha470, 16'ha450, 16'h9c50, 16'h9c4f, 16'h9c4f, 16'h93ee, 16'h4a6, 16'h293, 16'h212, 16'h212, 16'h20e2, 16'h18c1, 16'h820, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h6ac9, 16'h6ae9, 16'h6aea, 16'h73a, 16'h732a, 16'h734b, 16'h7b6b, 16'h836c, 16'h838c, 16'h83ad, 16'h8bad, 16'h8bcd, 16'h8bed, 16'h8bed, 16'h8bee, 16'h94e, 16'h94e, 16'h8bed, 16'h39c5, 16'h881, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h881, 16'h2986, 16'h4a28, 16'h18c2, 16'h1081, 16'h020, 16'h020, 16'h020, 16'h020, 16'h040, 16'h040, 16'h040, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h1061, 16'h6268, 16'h72c9, 16'h6ac9, 16'h6ac9, 16'h6ac9, 16'h4a6, 16'h3964, 16'h3144, 16'h2923, 16'h213, 16'h213, 16'h20e3, 16'h213, 16'h20e3, 16'h18c2, 16'h20e3, 16'h18e2, 16'h20e2, 16'h294, 16'h7b6c, 16'h6bb, 16'h2948, 16'h298c, 16'h10c9, 16'h887, 16'h5a6b, 16'h8bab, 16'h5a47, 16'h5227, 16'h5247, 16'h5a47, 16'h5a47, 16'h5a47, 16'h5a47, 16'h5a47, 16'h5a68, 16'h6288, 16'h72c9, 16'h93ed, 16'h6ac9, 16'h41c5, 16'h1081, 16'h820, 16'h820, 16'h820, 16'h820, 16'h820, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h820, 16'h840, 16'h840, 16'h840, 16'h840, 16'h3965, 16'hacb1, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha470, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha450, 16'ha450, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'ha44f, 16'ha470, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h93ee, 16'h4a6, 16'h213, 16'h212, 16'h20e2, 16'h20e2, 16'h18c1, 16'h820, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h62a9, 16'h62a9, 16'h6ac9, 16'h6ae9, 16'h6aea, 16'h73a, 16'h732b, 16'h732b, 16'h7b6c, 16'h7b6c, 16'h838c, 16'h83ac, 16'h83ad, 16'h8bcd, 16'h8bcd, 16'h8bed, 16'h8bed, 16'h83cd, 16'h39c5, 16'h881, 16'h060, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h1081, 16'h2985, 16'h4a47, 16'h18e2, 16'h1081, 16'h020, 16'h020, 16'h020, 16'h040, 16'h040, 16'h040, 16'h040, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h1061, 16'h6268, 16'h72e9, 16'h72c9, 16'h72c9, 16'h6aa9, 16'h49c6, 16'h3144, 16'h2944, 16'h2923, 16'h213, 16'h213, 16'h20e3, 16'h20e3, 16'h213, 16'h213, 16'h18a2, 16'h20e2, 16'h20e2, 16'h20e3, 16'h427, 16'h4a28, 16'h2948, 16'h296c, 16'h10e9, 16'h887, 16'h2947, 16'h72e8, 16'h6287, 16'h5a47, 16'h5a47, 16'h5a47, 16'h5a47, 16'h5a47, 16'h5a47, 16'h5a47, 16'h5a67, 16'h6288, 16'h72c9, 16'h93ed, 16'h6ac9, 16'h41c5, 16'h1061, 16'h020, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h820, 16'h840, 16'h840, 16'h840, 16'h3965, 16'hacb1, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha470, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha46f, 16'ha46f, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h93ed, 16'h4a6, 16'h212, 16'h212, 16'h212, 16'h20e2, 16'h18c1, 16'h820, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h6288, 16'h62a9, 16'h62a9, 16'h62c9, 16'h6ac9, 16'h6ae9, 16'h6aea, 16'h73a, 16'h732b, 16'h7b4b, 16'h7b6b, 16'h7b6c, 16'h838c, 16'h83ac, 16'h83ac, 16'h8bcd, 16'h8bcd, 16'h83ac, 16'h39a4, 16'h880, 16'h060, 16'h060, 16'h860, 16'h860, 16'h840, 16'h040, 16'h1081, 16'h2985, 16'h4a47, 16'h18c2, 16'h1061, 16'h020, 16'h020, 16'h020, 16'h020, 16'h040, 16'h040, 16'h040, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h00, 16'h020, 16'h840, 16'h840, 16'h020, 16'h020, 16'h1081, 16'h6288, 16'h72c9, 16'h6ac9, 16'h72c9, 16'h62a8, 16'h41c6, 16'h3164, 16'h2944, 16'h2123, 16'h213, 16'h20e3, 16'h20e2, 16'h20e2, 16'h18e2, 16'h213, 16'h1082, 16'h10a1, 16'h20e2, 16'h20e2, 16'h18e2, 16'h20e3, 16'h2926, 16'h298b, 16'h199, 16'h10a7, 16'h4a9, 16'h7b8, 16'h6287, 16'h5a47, 16'h5a47, 16'h5a47, 16'h5a47, 16'h5a47, 16'h5a47, 16'h5a67, 16'h5a67, 16'h6288, 16'h72e9, 16'h93ed, 16'h6ac9, 16'h41c5, 16'h1061, 16'h020, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h840, 16'h840, 16'h3164, 16'hacb1, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb0, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'hac90, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha46f, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'ha44f, 16'ha46f, 16'ha470, 16'ha470, 16'h9c70, 16'h9c4f, 16'h9c4f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h8bed, 16'h4a7, 16'h213, 16'h212, 16'h212, 16'h20e1, 16'h18c1, 16'h820, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h5a88, 16'h5a88, 16'h62a8, 16'h62a9, 16'h62c9, 16'h6ac9, 16'h62e9, 16'h6aea, 16'h73a, 16'h73a, 16'h732b, 16'h7b4b, 16'h7b6b, 16'h7b6c, 16'h838c, 16'h83ac, 16'h83ad, 16'h838c, 16'h39a4, 16'h860, 16'h860, 16'h860, 16'h860, 16'h860, 16'h860, 16'h861, 16'h18e2, 16'h39c7, 16'h4a48, 16'h18c2, 16'h1061, 16'h020, 16'h020, 16'h020, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h1081, 16'h41c5, 16'h2944, 16'h840, 16'h020, 16'h1881, 16'h6288, 16'h72c9, 16'h72e9, 16'h72c9, 16'h6288, 16'h39a5, 16'h3164, 16'h2924, 16'h2923, 16'h293, 16'h20e2, 16'h20e2, 16'h20e2, 16'h18e2, 16'h20e3, 16'h18e3, 16'h18a2, 16'h1081, 16'h20e2, 16'h20e3, 16'h3165, 16'h41c7, 16'h2969, 16'h192a, 16'h10c8, 16'h5229, 16'h7ae8, 16'h6287, 16'h5a67, 16'h5a67, 16'h5a47, 16'h5a47, 16'h5a47, 16'h5a47, 16'h5a67, 16'h5a67, 16'h6288, 16'h72c9, 16'h93ed, 16'h6ac9, 16'h41c5, 16'h1061, 16'h020, 16'h820, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h840, 16'h840, 16'h3144, 16'hac90, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'hac90, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'ha44f, 16'ha46f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h8bed, 16'h4a6, 16'h212, 16'h212, 16'h20e2, 16'h20e2, 16'h18c1, 16'h840, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h5a68, 16'h5a88, 16'h5a88, 16'h62a8, 16'h62a9, 16'h62c9, 16'h62c9, 16'h6ac9, 16'h6ae9, 16'h6b9, 16'h6ba, 16'h732b, 16'h732b, 16'h7b4b, 16'h7b6b, 16'h7b8c, 16'h838c, 16'h7b6c, 16'h3184, 16'h1081, 16'h10a1, 16'h18c1, 16'h212, 16'h2923, 16'h3184, 16'h39a5, 16'h5247, 16'h62ea, 16'h5248, 16'h18c2, 16'h1061, 16'h020, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h00, 16'h20e3, 16'h62a8, 16'h39a5, 16'h840, 16'h020, 16'h1881, 16'h6288, 16'h72c9, 16'h72c9, 16'h6ac9, 16'h6288, 16'h3985, 16'h3144, 16'h2924, 16'h213, 16'h213, 16'h213, 16'h20c3, 16'h20e3, 16'h20e2, 16'h20e2, 16'h18e3, 16'h213, 16'h18c2, 16'h18a2, 16'h20e3, 16'h427, 16'h5aab, 16'h2968, 16'h214a, 16'h18c8, 16'h49c8, 16'h7b8, 16'h6287, 16'h5a67, 16'h5a47, 16'h5a47, 16'h5a47, 16'h5a47, 16'h5a47, 16'h5a67, 16'h5a67, 16'h6288, 16'h72c9, 16'h93ed, 16'h6ac9, 16'h41c5, 16'h861, 16'h020, 16'h820, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h820, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h040, 16'h840, 16'h3144, 16'hac90, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha46f, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2f, 16'h8bcd, 16'h4a6, 16'h213, 16'h212, 16'h20e2, 16'h20e2, 16'h18c2, 16'h820, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h5a68, 16'h5a68, 16'h5a88, 16'h62a8, 16'h62a8, 16'h62a9, 16'h62c9, 16'h62c9, 16'h6ac9, 16'h6ae9, 16'h6ae9, 16'h6ba, 16'h732a, 16'h734b, 16'h7b4b, 16'h7b6b, 16'h838b, 16'h7b8b, 16'h5a87, 16'h4a47, 16'h5aa8, 16'h6b9, 16'h734b, 16'h7b8c, 16'h83cd, 16'h8bcd, 16'h8bed, 16'h7b6c, 16'h5248, 16'h20e2, 16'h1061, 16'h020, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h00, 16'h18e3, 16'h5a88, 16'h3184, 16'h840, 16'h020, 16'h1881, 16'h6288, 16'h72c9, 16'h72ca, 16'h6ac9, 16'h5a88, 16'h39a5, 16'h3144, 16'h2923, 16'h293, 16'h213, 16'h20e3, 16'h20e3, 16'h20e3, 16'h18e2, 16'h20e2, 16'h18e3, 16'h18e3, 16'h213, 16'h3144, 16'h2924, 16'h39c6, 16'h5a8b, 16'h3145, 16'h3167, 16'h20e5, 16'h28e3, 16'h72a7, 16'h6287, 16'h5a47, 16'h5a67, 16'h5a47, 16'h5a67, 16'h5a67, 16'h5a67, 16'h5a67, 16'h5a67, 16'h6288, 16'h72c9, 16'h93ed, 16'h6ac9, 16'h41c5, 16'h861, 16'h020, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h820, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h840, 16'h3144, 16'hac90, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'ha4b0, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha44f, 16'h9c4f, 16'ha44f, 16'h9c4f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9ce, 16'h8bcd, 16'h4a7, 16'h213, 16'h212, 16'h20e2, 16'h20e2, 16'h18c1, 16'h820, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h5267, 16'h5a88, 16'h5a88, 16'h5a88, 16'h62a8, 16'h62a8, 16'h62a9, 16'h62a9, 16'h6ac9, 16'h6ae9, 16'h6ae9, 16'h6aea, 16'h6ba, 16'h732a, 16'h734a, 16'h7b4b, 16'h7b6b, 16'h838c, 16'h838c, 16'h83ac, 16'h83cd, 16'h8bed, 16'h8bed, 16'h8ce, 16'h94e, 16'h94e, 16'h944e, 16'h7b6c, 16'h5248, 16'h20e2, 16'h1061, 16'h020, 16'h040, 16'h040, 16'h040, 16'h040, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h00, 16'h00, 16'h841, 16'h18a2, 16'h861, 16'h020, 16'h020, 16'h1881, 16'h6288, 16'h72e9, 16'h72c9, 16'h6ac9, 16'h5a68, 16'h3985, 16'h3144, 16'h2923, 16'h213, 16'h213, 16'h20e3, 16'h20e2, 16'h20e2, 16'h18e2, 16'h18e2, 16'h18e2, 16'h20e2, 16'h18e2, 16'h3144, 16'h39a5, 16'h3184, 16'h41a6, 16'h3943, 16'h3984, 16'h3984, 16'h291, 16'h72c7, 16'h6287, 16'h5a67, 16'h5a67, 16'h5a47, 16'h5a67, 16'h5a67, 16'h5a67, 16'h5a67, 16'h5a67, 16'h6288, 16'h72c9, 16'h93ed, 16'h6ac9, 16'h41c5, 16'h861, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h840, 16'h840, 16'h3144, 16'hac90, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'ha4b0, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha44f, 16'ha44f, 16'ha46f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9ce, 16'h94e, 16'h8bcd, 16'h4a7, 16'h212, 16'h212, 16'h212, 16'h20e2, 16'h18c1, 16'h820, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h5267, 16'h5a67, 16'h5a88, 16'h5a88, 16'h6288, 16'h62a8, 16'h62a9, 16'h62a9, 16'h62c9, 16'h6ac9, 16'h6ae9, 16'h6ba, 16'h6ba, 16'h732a, 16'h734b, 16'h7b6b, 16'h838c, 16'h83ad, 16'h83cd, 16'h8bed, 16'h8ce, 16'h94e, 16'h942e, 16'h942f, 16'h942e, 16'h942f, 16'h9c4f, 16'h7b6c, 16'h5247, 16'h20e2, 16'h1061, 16'h020, 16'h040, 16'h020, 16'h020, 16'h040, 16'h040, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h1881, 16'h6288, 16'h72e9, 16'h6ac9, 16'h6ac9, 16'h6288, 16'h3985, 16'h3144, 16'h2944, 16'h2923, 16'h213, 16'h20e3, 16'h20e2, 16'h20e2, 16'h20e2, 16'h20e3, 16'h20e3, 16'h18c2, 16'h18e2, 16'h18c2, 16'h3164, 16'h41c5, 16'h59e4, 16'h6a42, 16'h59e2, 16'h41a3, 16'h3984, 16'h72e7, 16'h6a87, 16'h5a67, 16'h5a67, 16'h5a67, 16'h5a67, 16'h5a67, 16'h5a67, 16'h5a67, 16'h5a67, 16'h6288, 16'h72c9, 16'h93ed, 16'h6ac9, 16'h41c5, 16'h1061, 16'h020, 16'h00, 16'h020, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h840, 16'h840, 16'h3144, 16'ha490, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha46f, 16'ha470, 16'ha46f, 16'ha46f, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9ce, 16'h94e, 16'h8bcd, 16'h4a27, 16'h213, 16'h212, 16'h212, 16'h20e2, 16'h18c1, 16'h820, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h5267, 16'h5a68, 16'h5a88, 16'h5a88, 16'h62a9, 16'h62a9, 16'h62c9, 16'h6ac9, 16'h6ae9, 16'h6ba, 16'h6ba, 16'h732b, 16'h732b, 16'h734b, 16'h736b, 16'h736b, 16'h732b, 16'h838d, 16'h8bed, 16'h8ce, 16'h94e, 16'h94e, 16'h942f, 16'h94e, 16'h94e, 16'h8bed, 16'h83ad, 16'h73a, 16'h5268, 16'h20c2, 16'h861, 16'h020, 16'h040, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h1881, 16'h6a88, 16'h72c9, 16'h72c9, 16'h72c9, 16'h6288, 16'h39a5, 16'h3144, 16'h2924, 16'h213, 16'h213, 16'h213, 16'h213, 16'h20e3, 16'h18e3, 16'h18c3, 16'h18c3, 16'h18c2, 16'h18e2, 16'h18c2, 16'h20e2, 16'h6265, 16'ha3e5, 16'ha3e2, 16'h82e1, 16'h5a3, 16'h41a6, 16'h7ae9, 16'h6287, 16'h5a67, 16'h5a47, 16'h5a67, 16'h5a47, 16'h5a47, 16'h5a47, 16'h5a68, 16'h5a67, 16'h6287, 16'h6ac9, 16'h93ed, 16'h6ae9, 16'h49c5, 16'h1061, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h840, 16'h840, 16'h3144, 16'ha490, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha46f, 16'ha470, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h94e, 16'h94e, 16'h9ce, 16'h9ce, 16'h94e, 16'h8bcd, 16'h5226, 16'h213, 16'h212, 16'h212, 16'h20e2, 16'h18c1, 16'h840, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h5a68, 16'h5a88, 16'h5a88, 16'h5a88, 16'h5a89, 16'h5a89, 16'h5268, 16'h4a48, 16'h4a28, 16'h4a48, 16'h4a68, 16'h4a48, 16'h4a27, 16'h41e6, 16'h39c6, 16'h39a5, 16'h3165, 16'h62aa, 16'h8bee, 16'h8ce, 16'h734b, 16'h62ca, 16'h5268, 16'h41e6, 16'h3185, 16'h2124, 16'h18c2, 16'h20e3, 16'h41c6, 16'h20e2, 16'h1061, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h00, 16'h020, 16'h00, 16'h00, 16'h00, 16'h020, 16'h1881, 16'h6a88, 16'h72e9, 16'h72c9, 16'h72c9, 16'h6aa8, 16'h41a5, 16'h3144, 16'h2924, 16'h213, 16'h213, 16'h213, 16'h20e2, 16'h18e3, 16'h20e3, 16'h20e3, 16'h18e3, 16'h20c2, 16'h20e2, 16'h18c2, 16'h18c2, 16'h51c3, 16'h9bc4, 16'hb464, 16'h9bc4, 16'h5a5, 16'h49e8, 16'h8349, 16'h6287, 16'h5a67, 16'h5a47, 16'h5a47, 16'h5a67, 16'h5a67, 16'h5a67, 16'h5a67, 16'h5a67, 16'h6288, 16'h72c9, 16'h93ed, 16'h6ae9, 16'h49c5, 16'h1061, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h840, 16'h840, 16'h3144, 16'ha490, 16'hb4f1, 16'hb4f1, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4f1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb0, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'hacb0, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha46f, 16'ha470, 16'ha46f, 16'ha46f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9ce, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h8bcd, 16'h5227, 16'h212, 16'h212, 16'h211, 16'h20e2, 16'h18c1, 16'h840, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h3186, 16'h2965, 16'h2945, 16'h2125, 16'h2125, 16'h1926, 16'h2146, 16'h2125, 16'h2925, 16'h2945, 16'h2965, 16'h2124, 16'h2924, 16'h194, 16'h18e4, 16'h213, 16'h2124, 16'h5aa9, 16'h8ce, 16'h8bed, 16'h39a5, 16'h1081, 16'h840, 16'h040, 16'h040, 16'h040, 16'h040, 16'h1082, 16'h39a5, 16'h20c2, 16'h1061, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h1881, 16'h6aa8, 16'h6ac9, 16'h6ac9, 16'h6ac9, 16'h6aa9, 16'h41c6, 16'h3144, 16'h2923, 16'h213, 16'h213, 16'h20e3, 16'h20e2, 16'h18e3, 16'h20e3, 16'h20e3, 16'h18e2, 16'h18e2, 16'h18e2, 16'h20e2, 16'h20c2, 16'h20c2, 16'h49a4, 16'h9387, 16'h6a85, 16'h49e8, 16'h3987, 16'h6aa8, 16'h6287, 16'h5a47, 16'h5a47, 16'h5a67, 16'h5a67, 16'h5a67, 16'h5a67, 16'h5a67, 16'h6267, 16'h6288, 16'h72c9, 16'h93ed, 16'h72e9, 16'h49c5, 16'h1061, 16'h020, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h840, 16'h840, 16'h3124, 16'ha490, 16'hb4f1, 16'hb4f1, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha44f, 16'ha470, 16'ha46f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9ce, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h8bcd, 16'h5227, 16'h212, 16'h212, 16'h212, 16'h20e2, 16'h18c1, 16'h840, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h10c3, 16'h10c4, 16'h18e4, 16'h1925, 16'h2146, 16'h2986, 16'h39c7, 16'h39c6, 16'h41c7, 16'h39a7, 16'h3186, 16'h39a6, 16'h3165, 16'h2945, 16'h214, 16'h2924, 16'h2944, 16'h5269, 16'h94e, 16'h8cd, 16'h39a4, 16'h860, 16'h040, 16'h040, 16'h040, 16'h020, 16'h020, 16'h1082, 16'h3985, 16'h20c2, 16'h840, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h040, 16'h840, 16'h840, 16'h840, 16'h020, 16'h020, 16'h020, 16'h1881, 16'h6a88, 16'h6ac9, 16'h6ac9, 16'h6ac9, 16'h6aa9, 16'h49e6, 16'h3144, 16'h2923, 16'h2923, 16'h213, 16'h20e3, 16'h20e2, 16'h20c3, 16'h20e3, 16'h20e3, 16'h18e2, 16'h18e2, 16'h18e2, 16'h20e2, 16'h18c2, 16'h20e2, 16'h3965, 16'h93ed, 16'h72ea, 16'h41a7, 16'h20e6, 16'h72c8, 16'h6a87, 16'h5a47, 16'h5a47, 16'h5a67, 16'h5a47, 16'h5a67, 16'h5a67, 16'h5a67, 16'h6268, 16'h6288, 16'h72c9, 16'h93ed, 16'h72e9, 16'h49e5, 16'h1061, 16'h020, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h840, 16'h840, 16'h3124, 16'ha490, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f2, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb1, 16'hacb1, 16'hacb0, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha44f, 16'ha46f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h9c4e, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9ce, 16'h9c2e, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9ce, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h93ee, 16'h8bcd, 16'h5227, 16'h213, 16'h212, 16'h20e2, 16'h20e2, 16'h18c1, 16'h840, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h2124, 16'h2145, 16'h2965, 16'h3186, 16'h39c7, 16'h41e7, 16'h39a7, 16'h39c7, 16'h41e7, 16'h41e8, 16'h4a8, 16'h5269, 16'h41e7, 16'h3166, 16'h2125, 16'h2924, 16'h2965, 16'h4a8, 16'h8ce, 16'h942e, 16'h39c5, 16'h1081, 16'h040, 16'h020, 16'h020, 16'h020, 16'h020, 16'h1081, 16'h3184, 16'h18c2, 16'h820, 16'h840, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h040, 16'h840, 16'h861, 16'h1081, 16'h18a1, 16'h20e2, 16'h293, 16'h3164, 16'h3143, 16'h861, 16'h00, 16'h00, 16'h00, 16'h1882, 16'h6aa8, 16'h72c9, 16'h72c9, 16'h72c9, 16'h6ac8, 16'h5226, 16'h3164, 16'h2924, 16'h2123, 16'h213, 16'h20e3, 16'h20e3, 16'h20e3, 16'h20e3, 16'h20e2, 16'h20e3, 16'h18e3, 16'h18c2, 16'h18e2, 16'h18c2, 16'h18c2, 16'h3165, 16'h9c4e, 16'h9c4e, 16'h5a69, 16'h296, 16'h72c9, 16'h6a88, 16'h5a47, 16'h5a47, 16'h5a67, 16'h5a67, 16'h5a67, 16'h5a67, 16'h5a67, 16'h6267, 16'h6288, 16'h72c9, 16'h93ed, 16'h72e9, 16'h41e5, 16'h1061, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h840, 16'h3124, 16'ha470, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha46f, 16'ha470, 16'ha470, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9ce, 16'h9ce, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h93ee, 16'h8bad, 16'h5227, 16'h293, 16'h212, 16'h20e2, 16'h20e1, 16'h18c1, 16'h840, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h2945, 16'h2965, 16'h3186, 16'h39a6, 16'h39c7, 16'h41e7, 16'h39c7, 16'h39c7, 16'h39c7, 16'h41e7, 16'h41e7, 16'h41e8, 16'h39c8, 16'h3166, 16'h2925, 16'h2944, 16'h3165, 16'h41c6, 16'h8bee, 16'h944e, 16'h41c5, 16'h1081, 16'h040, 16'h020, 16'h020, 16'h020, 16'h020, 16'h1061, 16'h3164, 16'h1081, 16'h841, 16'h840, 16'h840, 16'h861, 16'h881, 16'h040, 16'h040, 16'h040, 16'h061, 16'h861, 16'h10a1, 16'h3964, 16'h41c5, 16'h41c5, 16'h49e6, 16'h4a6, 16'h5226, 16'h41c4, 16'h861, 16'h00, 16'h00, 16'h00, 16'h18a2, 16'h6aa8, 16'h6ac9, 16'h6ac9, 16'h6ac9, 16'h6ac8, 16'h5a67, 16'h3964, 16'h2924, 16'h2923, 16'h213, 16'h213, 16'h20e3, 16'h20e3, 16'h18e2, 16'h20e2, 16'h18e3, 16'h18e2, 16'h18e2, 16'h18e2, 16'h18c2, 16'h18c2, 16'h3165, 16'h9c4e, 16'ha46f, 16'ha46f, 16'h73c, 16'h7b9, 16'h6a88, 16'h5a48, 16'h5a47, 16'h5a67, 16'h5a67, 16'h5a67, 16'h5a67, 16'h5a68, 16'h6268, 16'h6288, 16'h72c9, 16'h93ed, 16'h72e9, 16'h41e5, 16'h1061, 16'h00, 16'h00, 16'h020, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h840, 16'h3124, 16'ha470, 16'hb4d2, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha450, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c2e, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h94e, 16'h94e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9ce, 16'h9ce, 16'h9ce, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h93ee, 16'h93ee, 16'h8bad, 16'h5227, 16'h293, 16'h212, 16'h212, 16'h20e2, 16'h18c1, 16'h840, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h2124, 16'h2125, 16'h2145, 16'h2125, 16'h2125, 16'h2145, 16'h2125, 16'h214, 16'h2125, 16'h2124, 16'h214, 16'h3186, 16'h39a7, 16'h39a7, 16'h3986, 16'h41e5, 16'h4a47, 16'h62a9, 16'h942f, 16'h9c6f, 16'h41e6, 16'h1081, 16'h040, 16'h020, 16'h020, 16'h020, 16'h020, 16'h841, 16'h18c2, 16'h840, 16'h861, 16'h10a2, 16'h2165, 16'h29a6, 16'h2165, 16'h881, 16'h061, 16'h061, 16'h881, 16'h881, 16'h881, 16'h3984, 16'h49e6, 16'h49e6, 16'h49e6, 16'h4a6, 16'h5226, 16'h41c4, 16'h861, 16'h00, 16'h00, 16'h00, 16'h18a2, 16'h6aa8, 16'h6ac9, 16'h6ac8, 16'h6ac8, 16'h6ac9, 16'h6288, 16'h39a5, 16'h2924, 16'h293, 16'h293, 16'h213, 16'h213, 16'h20e3, 16'h18e2, 16'h20e2, 16'h18e2, 16'h18e2, 16'h18e2, 16'h18c2, 16'h18c2, 16'h18c2, 16'h3165, 16'h9c4f, 16'ha490, 16'ha44f, 16'hb4f1, 16'ha42c, 16'h6aa8, 16'h5a68, 16'h5a47, 16'h5a48, 16'h5a68, 16'h5a68, 16'h5a67, 16'h5a68, 16'h6268, 16'h6288, 16'h72e9, 16'h94d, 16'h72e9, 16'h41e5, 16'h1061, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h820, 16'h840, 16'h3124, 16'ha470, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'ha490, 16'ha490, 16'ha470, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha450, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c4f, 16'h9c4f, 16'h9c4e, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h94e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2f, 16'h9c2e, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9ce, 16'h9ce, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h93ee, 16'h93ed, 16'h8bcd, 16'h5227, 16'h293, 16'h212, 16'h212, 16'h20e2, 16'h18c1, 16'h840, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h18c3, 16'h18e4, 16'h214, 16'h215, 16'h2125, 16'h2965, 16'h3186, 16'h39c6, 16'h4a27, 16'h5248, 16'h5aa9, 16'h6bb, 16'h7b4b, 16'h7b8c, 16'h83cd, 16'h94d, 16'h9c4f, 16'h9c70, 16'ha4b1, 16'ha490, 16'h41e6, 16'h1081, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h10a2, 16'h1924, 16'h29a6, 16'h31e7, 16'h2186, 16'h881, 16'h061, 16'h061, 16'h881, 16'h061, 16'h881, 16'h3984, 16'h49e5, 16'h49e6, 16'h49e6, 16'h49e6, 16'h526, 16'h41c4, 16'h841, 16'h00, 16'h00, 16'h00, 16'h18a2, 16'h6aa8, 16'h6ac9, 16'h6ac9, 16'h6ac9, 16'h6ac9, 16'h6aa8, 16'h49e6, 16'h3144, 16'h2923, 16'h2923, 16'h213, 16'h20e3, 16'h20e3, 16'h20e2, 16'h20e2, 16'h20e3, 16'h18e2, 16'h18c2, 16'h18c2, 16'h18c2, 16'h20c2, 16'h3185, 16'h9c4f, 16'hacb0, 16'ha42f, 16'hb4f1, 16'hac6d, 16'h6aa8, 16'h5a68, 16'h5a47, 16'h5a47, 16'h5a67, 16'h5a67, 16'h5a67, 16'h5a68, 16'h6268, 16'h6288, 16'h72e9, 16'h94d, 16'h72e9, 16'h41c5, 16'h1061, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h840, 16'h3124, 16'ha470, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha470, 16'ha46f, 16'ha470, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9ce, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94d, 16'h93ed, 16'h8bcd, 16'h5227, 16'h293, 16'h212, 16'h20e2, 16'h20e2, 16'h18c1, 16'h840, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h4a26, 16'h5268, 16'h62a9, 16'h6ba, 16'h734a, 16'h7b6b, 16'h838c, 16'h8bcc, 16'h8bed, 16'h8cd, 16'h94e, 16'h94e, 16'h942f, 16'h9c4f, 16'h9c6f, 16'ha490, 16'ha490, 16'ha4b1, 16'hacd1, 16'ha4b0, 16'h41e6, 16'h1081, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h861, 16'h10c3, 16'h2186, 16'h29c7, 16'h2165, 16'h861, 16'h061, 16'h061, 16'h061, 16'h060, 16'h860, 16'h3984, 16'h49e5, 16'h49e5, 16'h49e6, 16'h49e6, 16'h526, 16'h41a4, 16'h841, 16'h00, 16'h00, 16'h00, 16'h18a2, 16'h6aa8, 16'h6ac9, 16'h6ac9, 16'h6ac9, 16'h6ac9, 16'h6ac9, 16'h5247, 16'h3164, 16'h2923, 16'h2923, 16'h213, 16'h213, 16'h213, 16'h20e2, 16'h20e3, 16'h18c3, 16'h18c2, 16'h18c2, 16'h18e3, 16'h20c2, 16'h18c2, 16'h3185, 16'h9c6f, 16'hb4f1, 16'ha44f, 16'ha46f, 16'hac6d, 16'h6aa7, 16'h5a68, 16'h5a47, 16'h5a67, 16'h5a47, 16'h5a67, 16'h5a67, 16'h5a68, 16'h6268, 16'h6288, 16'h72e9, 16'h94d, 16'h72e9, 16'h41c5, 16'h1061, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h840, 16'h2924, 16'ha470, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha46f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9ce, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9ce, 16'h9ce, 16'h9ce, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h93ee, 16'h94e, 16'h93ee, 16'h93ee, 16'h93ee, 16'h8bad, 16'h5227, 16'h213, 16'h20e2, 16'h20e2, 16'h20e2, 16'h18c2, 16'h840, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h7b6b, 16'h838b, 16'h83ac, 16'h8bcc, 16'h8bcc, 16'h8bed, 16'h8bed, 16'h93ed, 16'h94e, 16'h94e, 16'h942e, 16'h942f, 16'h944e, 16'h9c4e, 16'h9c6f, 16'ha490, 16'ha4b0, 16'hacd1, 16'hacd1, 16'ha4b0, 16'h49e6, 16'h1081, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h00, 16'h10a2, 16'h2186, 16'h29a6, 16'h2165, 16'h061, 16'h060, 16'h060, 16'h060, 16'h040, 16'h861, 16'h3964, 16'h41c5, 16'h49e5, 16'h49e5, 16'h49e5, 16'h4a6, 16'h39a4, 16'h841, 16'h00, 16'h00, 16'h00, 16'h1882, 16'h6aa8, 16'h6ac9, 16'h6ac9, 16'h6ac9, 16'h6ac9, 16'h6ac9, 16'h6aa9, 16'h41c5, 16'h3123, 16'h293, 16'h213, 16'h213, 16'h20e3, 16'h20e3, 16'h20e3, 16'h18c3, 16'h20e3, 16'h20c2, 16'h18e2, 16'h18c2, 16'h18c2, 16'h3985, 16'h9c6f, 16'hb4d1, 16'hacd1, 16'ha44e, 16'ha44c, 16'h6aa8, 16'h5a67, 16'h5a67, 16'h5a67, 16'h5a67, 16'h5a67, 16'h5a67, 16'h5a68, 16'h6268, 16'h6288, 16'h72e9, 16'h94d, 16'h72e9, 16'h41c5, 16'h1061, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h840, 16'h2924, 16'ha46f, 16'hb4d1, 16'hb4f1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha46f, 16'ha44f, 16'h9c4f, 16'h9c50, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9ce, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9cf, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2f, 16'h9c2f, 16'h9ce, 16'h9ce, 16'h9ce, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h93ed, 16'h93ed, 16'h93ee, 16'h93ee, 16'h93ed, 16'h8bad, 16'h5227, 16'h213, 16'h212, 16'h20e2, 16'h20e2, 16'h18c1, 16'h840, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h838b, 16'h83ac, 16'h8bac, 16'h8bcc, 16'h8bed, 16'h8bed, 16'h93ed, 16'h94d, 16'h94e, 16'h94e, 16'h942e, 16'h942e, 16'h944e, 16'h9c4f, 16'h9c6f, 16'ha490, 16'ha4b0, 16'hacd1, 16'hacf1, 16'ha4b0, 16'h41e6, 16'h1081, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h00, 16'h10a2, 16'h2185, 16'h21a6, 16'h2165, 16'h061, 16'h060, 16'h060, 16'h060, 16'h060, 16'h861, 16'h3964, 16'h41c5, 16'h41c5, 16'h49c5, 16'h49e5, 16'h4a5, 16'h3984, 16'h841, 16'h00, 16'h00, 16'h00, 16'h18a2, 16'h6aa8, 16'h6ac9, 16'h6ac9, 16'h6ac9, 16'h6ac9, 16'h6aa9, 16'h72c9, 16'h6aa8, 16'h41c5, 16'h293, 16'h213, 16'h213, 16'h213, 16'h20e3, 16'h20e3, 16'h18e3, 16'h20e3, 16'h20e2, 16'h18e2, 16'h20e2, 16'h20e2, 16'h3965, 16'ha44f, 16'hb4f1, 16'hb4f1, 16'hac8f, 16'ha4b, 16'h6aa8, 16'h6267, 16'h5a67, 16'h5a67, 16'h5a68, 16'h5a67, 16'h5a67, 16'h5a67, 16'h6267, 16'h6288, 16'h72e9, 16'h94d, 16'h72e9, 16'h41e5, 16'h861, 16'h00, 16'h00, 16'h00, 16'h020, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h840, 16'h2924, 16'ha46f, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha46f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2f, 16'h9c2e, 16'h94e, 16'h94e, 16'h9ce, 16'h9c2e, 16'h9c2e, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9ce, 16'h9ce, 16'h9c2f, 16'h9ce, 16'h9ce, 16'h9ce, 16'h9ce, 16'h94e, 16'h93ee, 16'h94e, 16'h94e, 16'h94d, 16'h93ee, 16'h93ee, 16'h93ed, 16'h93ed, 16'h93ed, 16'h8bad, 16'h5227, 16'h293, 16'h212, 16'h20e2, 16'h20e2, 16'h18c1, 16'h840, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h838b, 16'h83ac, 16'h8bcc, 16'h8bec, 16'h8bed, 16'h8bed, 16'h94d, 16'h94d, 16'h94d, 16'h942e, 16'h942e, 16'h942e, 16'h9c4f, 16'h9c4f, 16'h9c6f, 16'ha490, 16'ha4b0, 16'hacd1, 16'hacd1, 16'ha4b0, 16'h41e5, 16'h1081, 16'h040, 16'h020, 16'h040, 16'h040, 16'h020, 16'h020, 16'h020, 16'h020, 16'h00, 16'h882, 16'h2165, 16'h29a6, 16'h2985, 16'h061, 16'h060, 16'h861, 16'h881, 16'h881, 16'h1081, 16'h3984, 16'h41c5, 16'h41c5, 16'h41c5, 16'h49c5, 16'h49e5, 16'h3984, 16'h841, 16'h00, 16'h00, 16'h00, 16'h293, 16'h72c9, 16'h6aa9, 16'h6ac9, 16'h6aa9, 16'h6ac9, 16'h6ac8, 16'h72c9, 16'h7b2a, 16'h6287, 16'h2924, 16'h20e3, 16'h213, 16'h213, 16'h213, 16'h20e3, 16'h20e3, 16'h20e3, 16'h20e3, 16'h20e3, 16'h20e2, 16'h20e2, 16'h3985, 16'h9c6f, 16'hb4f1, 16'hb4f1, 16'hb511, 16'hac6d, 16'h6aa8, 16'h5a67, 16'h5a67, 16'h5a67, 16'h5a68, 16'h5a67, 16'h5a68, 16'h5a68, 16'h6267, 16'h62a8, 16'h72e9, 16'h94d, 16'h6ae9, 16'h41c5, 16'h861, 16'h020, 16'h00, 16'h00, 16'h020, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h840, 16'h840, 16'h2924, 16'ha46f, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacd1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9ce, 16'h9ce, 16'h9ce, 16'h9ce, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9ce, 16'h9ce, 16'h9ce, 16'h94e, 16'h94e, 16'h94e, 16'h93ee, 16'h93ee, 16'h93ed, 16'h94e, 16'h93ee, 16'h93ee, 16'h93ed, 16'h93ed, 16'h93ed, 16'h8bac, 16'h5227, 16'h293, 16'h212, 16'h20e2, 16'h20e1, 16'h18c1, 16'h840, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h838b, 16'h83ac, 16'h8bcd, 16'h8bcd, 16'h8bed, 16'h8bed, 16'h93ed, 16'h94d, 16'h94d, 16'h942e, 16'h942e, 16'h942f, 16'h944e, 16'h9c4f, 16'h9c6f, 16'ha490, 16'ha490, 16'ha4b0, 16'hacd1, 16'ha490, 16'h41e5, 16'h1081, 16'h040, 16'h020, 16'h040, 16'h040, 16'h020, 16'h020, 16'h020, 16'h020, 16'h00, 16'h041, 16'h10c2, 16'h113, 16'h2164, 16'h18e2, 16'h213, 16'h3164, 16'h41e5, 16'h3163, 16'h18a1, 16'h41a4, 16'h41c5, 16'h41c5, 16'h41c5, 16'h41c5, 16'h49e5, 16'h3983, 16'h840, 16'h00, 16'h00, 16'h00, 16'h28e3, 16'h6aa9, 16'h6aa9, 16'h6aa9, 16'h6aa9, 16'h6aa9, 16'h6aa9, 16'h72c9, 16'h7b2a, 16'h62a8, 16'h20e2, 16'h861, 16'h10a2, 16'h18c2, 16'h20e2, 16'h20e3, 16'h18e3, 16'h20e3, 16'h20e3, 16'h20e3, 16'h20e2, 16'h20c2, 16'h3985, 16'ha46f, 16'hb4f1, 16'hb511, 16'hb511, 16'hac6d, 16'h6aa8, 16'h5a67, 16'h5a67, 16'h5a67, 16'h5a67, 16'h5a67, 16'h5a68, 16'h5a68, 16'h6268, 16'h6288, 16'h72e9, 16'h94d, 16'h6ae9, 16'h41c5, 16'h1061, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h840, 16'h840, 16'h2924, 16'ha46f, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'ha490, 16'ha470, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha46f, 16'ha44f, 16'ha46f, 16'ha470, 16'ha46f, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9ce, 16'h94e, 16'h9ce, 16'h9ce, 16'h94e, 16'h9ce, 16'h9c2e, 16'h9ce, 16'h9ce, 16'h9ce, 16'h9c2e, 16'h9ce, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94d, 16'h93ed, 16'h93ed, 16'h93ee, 16'h93ee, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h8bac, 16'h5227, 16'h292, 16'h212, 16'h20e2, 16'h20e2, 16'h20c1, 16'h840, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h838b, 16'h83ac, 16'h8bcc, 16'h8bcd, 16'h8bcd, 16'h8bed, 16'h8bed, 16'h93ed, 16'h94d, 16'h94e, 16'h94e, 16'h942e, 16'h942e, 16'h9c4f, 16'h9c4f, 16'h9c6f, 16'ha490, 16'ha4b0, 16'ha4b0, 16'ha48f, 16'h41e6, 16'h1061, 16'h040, 16'h040, 16'h040, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h861, 16'h18a1, 16'h841, 16'h3144, 16'h49e5, 16'h4a6, 16'h4a6, 16'h5a67, 16'h3984, 16'h840, 16'h3963, 16'h41a5, 16'h41a5, 16'h41a4, 16'h41c5, 16'h49e5, 16'h3983, 16'h840, 16'h00, 16'h00, 16'h00, 16'h28e3, 16'h6aa8, 16'h6aa9, 16'h6aa9, 16'h6aa9, 16'h6aa8, 16'h6aa9, 16'h6ac9, 16'h7b2a, 16'h62a8, 16'h20c2, 16'h020, 16'h020, 16'h820, 16'h841, 16'h1061, 16'h10a2, 16'h18a2, 16'h18c2, 16'h18c2, 16'h18c2, 16'h18c2, 16'h3986, 16'ha470, 16'hb512, 16'hbd12, 16'hbd11, 16'hac6d, 16'h6a88, 16'h5a47, 16'h5a67, 16'h5a47, 16'h5a67, 16'h5a67, 16'h5a67, 16'h5a67, 16'h6268, 16'h6288, 16'h72e9, 16'h94d, 16'h72e9, 16'h41c5, 16'h1061, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h840, 16'h2924, 16'ha46f, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha470, 16'ha46f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9ce, 16'h9ce, 16'h94e, 16'h9ce, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h9ce, 16'h9ce, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ee, 16'h93ee, 16'h93ed, 16'h93ed, 16'h93cd, 16'h93cd, 16'h8bac, 16'h5227, 16'h292, 16'h212, 16'h20e2, 16'h20e2, 16'h18c1, 16'h840, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h838b, 16'h83ac, 16'h8bac, 16'h8bcc, 16'h8bcc, 16'h8bcd, 16'h8bed, 16'h8bed, 16'h93ed, 16'h94d, 16'h94e, 16'h94e, 16'h94e, 16'h942f, 16'h9c4f, 16'h9c4f, 16'h9c70, 16'ha490, 16'ha4b0, 16'h9c6f, 16'h41e5, 16'h1081, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h020, 16'h020, 16'h020, 16'h020, 16'h1081, 16'h18e2, 16'h840, 16'h3144, 16'h4a6, 16'h526, 16'h526, 16'h5a67, 16'h3984, 16'h840, 16'h3963, 16'h41a4, 16'h41a5, 16'h41a5, 16'h41a5, 16'h49c5, 16'h3964, 16'h840, 16'h00, 16'h841, 16'h18a2, 16'h3984, 16'h72a8, 16'h6aa8, 16'h6aa9, 16'h6aa9, 16'h6aa9, 16'h6aa9, 16'h6ac9, 16'h7b2a, 16'h6aa8, 16'h20c2, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h020, 16'h820, 16'h820, 16'h841, 16'h861, 16'h3145, 16'ha490, 16'hbd12, 16'hbd32, 16'hb4f1, 16'ha42c, 16'h6a88, 16'h5a67, 16'h5a67, 16'h5a67, 16'h5a67, 16'h5a67, 16'h5a67, 16'h5a68, 16'h6268, 16'h6288, 16'h72e9, 16'h94d, 16'h72e9, 16'h41c5, 16'h861, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h840, 16'h2924, 16'ha46f, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha44f, 16'ha46f, 16'ha470, 16'ha470, 16'ha470, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h94e, 16'h9ce, 16'h9c2e, 16'h9c2e, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h93ee, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93cd, 16'h93cd, 16'h8bac, 16'h5247, 16'h212, 16'h212, 16'h20e2, 16'h20e2, 16'h18c1, 16'h840, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h836b, 16'h838c, 16'h83ac, 16'h8bac, 16'h8bcc, 16'h8bcd, 16'h8bcd, 16'h8bed, 16'h8bed, 16'h8bed, 16'h94d, 16'h94e, 16'h94e, 16'h942e, 16'h942f, 16'h9c4f, 16'h9c6f, 16'h9c70, 16'ha490, 16'h9c4f, 16'h41c5, 16'h1061, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h840, 16'h020, 16'h3144, 16'h4a6, 16'h4a7, 16'h5226, 16'h5a67, 16'h3984, 16'h841, 16'h3963, 16'h41a4, 16'h41a5, 16'h41a5, 16'h41a5, 16'h49c5, 16'h3964, 16'h840, 16'h820, 16'h18a2, 16'h841, 16'h20c2, 16'h6a88, 16'h6aa9, 16'h6aa9, 16'h6aa9, 16'h6aa8, 16'h6aa9, 16'h6ac9, 16'h7b2a, 16'h6288, 16'h20c2, 16'h020, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h2924, 16'ha490, 16'hbd12, 16'hb511, 16'h93ed, 16'h8b69, 16'h6a88, 16'h5a67, 16'h5a67, 16'h5a67, 16'h5a67, 16'h5a67, 16'h5a67, 16'h6268, 16'h6288, 16'h6a88, 16'h72e9, 16'h9cd, 16'h72e9, 16'h41c5, 16'h861, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h840, 16'h840, 16'h2924, 16'ha46f, 16'hb4d1, 16'hb4d2, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha46f, 16'ha470, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9ce, 16'h9ce, 16'h9ce, 16'h9ce, 16'h9ce, 16'h9ce, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93cd, 16'h93cd, 16'h8bad, 16'h5247, 16'h212, 16'h212, 16'h20e2, 16'h20e2, 16'h20c1, 16'h840, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h7b6b, 16'h836c, 16'h838c, 16'h838c, 16'h83ac, 16'h83ac, 16'h8bad, 16'h8bcd, 16'h8bcd, 16'h8bed, 16'h8bed, 16'h8bed, 16'h94e, 16'h94e, 16'h94e, 16'h942e, 16'h9c4f, 16'h9c4f, 16'h9c6f, 16'h944e, 16'h41c5, 16'h1060, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h020, 16'h00, 16'h020, 16'h820, 16'h3164, 16'h4a26, 16'h5226, 16'h5226, 16'h5a67, 16'h3984, 16'h841, 16'h3963, 16'h41a5, 16'h41a5, 16'h41a4, 16'h41a4, 16'h41c5, 16'h3163, 16'h840, 16'h1061, 16'h20e3, 16'h00, 16'h1882, 16'h6288, 16'h6aa9, 16'h6aa8, 16'h6aa8, 16'h6aa8, 16'h6aa8, 16'h6ac9, 16'h7ba, 16'h6288, 16'h20c2, 16'h820, 16'h820, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h820, 16'h2924, 16'ha470, 16'hacb0, 16'hacb0, 16'h836b, 16'h8b69, 16'h6a87, 16'h5a67, 16'h5a67, 16'h5a67, 16'h5a67, 16'h5a67, 16'h5a67, 16'h6268, 16'h6268, 16'h6288, 16'h72e9, 16'h9c2d, 16'h72e9, 16'h41c4, 16'h861, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h840, 16'h840, 16'h3124, 16'ha46f, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'hac90, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha470, 16'ha46f, 16'ha44f, 16'ha44f, 16'ha470, 16'ha46f, 16'ha470, 16'ha46f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9ce, 16'h9ce, 16'h9ce, 16'h9ce, 16'h94e, 16'h94e, 16'h94e, 16'h9ce, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h93ee, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93cd, 16'h93cd, 16'h8bac, 16'h5227, 16'h212, 16'h212, 16'h20e2, 16'h20e2, 16'h18c1, 16'h840, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h7b6b, 16'h836b, 16'h836c, 16'h7b6b, 16'h836c, 16'h83ad, 16'h83ac, 16'h83ac, 16'h8bcc, 16'h8bcd, 16'h8bed, 16'h8bed, 16'h8bed, 16'h93ed, 16'h94e, 16'h942e, 16'h942f, 16'h9c2f, 16'h9c4f, 16'h942e, 16'h41c5, 16'h1080, 16'h040, 16'h860, 16'h040, 16'h060, 16'h060, 16'h040, 16'h040, 16'h840, 16'h840, 16'h040, 16'h040, 16'h840, 16'h3164, 16'h5226, 16'h5226, 16'h5226, 16'h5a67, 16'h3984, 16'h841, 16'h3963, 16'h41a4, 16'h41a4, 16'h41a4, 16'h41a4, 16'h41c5, 16'h3163, 16'h840, 16'h841, 16'h213, 16'h821, 16'h1882, 16'h6288, 16'h6aa9, 16'h6aa8, 16'h6aa9, 16'h62a8, 16'h6aa8, 16'h6ac9, 16'h7ba, 16'h6288, 16'h20c2, 16'h020, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h820, 16'h840, 16'h840, 16'h861, 16'h3124, 16'h9c2f, 16'ha44f, 16'h9c2e, 16'h72ea, 16'h8328, 16'h6a87, 16'h5a48, 16'h5a67, 16'h5a67, 16'h5a48, 16'h5a48, 16'h5a67, 16'h6267, 16'h6268, 16'h6288, 16'h72e9, 16'h9c2d, 16'h72e9, 16'h49e5, 16'h1061, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h840, 16'h840, 16'h2924, 16'h9c6f, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'ha490, 16'hac90, 16'hac90, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha450, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha46f, 16'ha46f, 16'ha470, 16'ha46f, 16'ha44f, 16'h9c4f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9ce, 16'h9ce, 16'h9ce, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94d, 16'h94d, 16'h93ee, 16'h93ee, 16'h94e, 16'h94d, 16'h94d, 16'h93ee, 16'h93ee, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93cd, 16'h93ed, 16'h93cd, 16'h93cd, 16'h8bcd, 16'h8bac, 16'h5227, 16'h293, 16'h20e2, 16'h20e2, 16'h20e2, 16'h18a1, 16'h840, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h732a, 16'h7b2b, 16'h7b2b, 16'h732a, 16'h7b2b, 16'h838c, 16'h838c, 16'h83ac, 16'h8bac, 16'h8bac, 16'h8bcd, 16'h8bcd, 16'h8bcd, 16'h8bed, 16'h8cd, 16'h94e, 16'h942f, 16'h942f, 16'h9c2f, 16'h94e, 16'h41c5, 16'h880, 16'h860, 16'h880, 16'h880, 16'h880, 16'h1080, 16'h1081, 16'h10c1, 16'h212, 16'h2944, 16'h18c2, 16'h861, 16'h840, 16'h3164, 16'h5226, 16'h5226, 16'h4a27, 16'h5a67, 16'h3984, 16'h840, 16'h3163, 16'h41a4, 16'h39a4, 16'h41a4, 16'h41a4, 16'h41c4, 16'h3143, 16'h820, 16'h00, 16'h18c3, 16'h213, 16'h18a2, 16'h6268, 16'h6aa8, 16'h6aa8, 16'h62a8, 16'h62a8, 16'h6289, 16'h6288, 16'h6aa9, 16'h4a26, 16'h18c2, 16'h020, 16'h020, 16'h020, 16'h040, 16'h040, 16'h040, 16'h840, 16'h840, 16'h860, 16'h860, 16'h1081, 16'h3144, 16'h9c2f, 16'h9c4f, 16'ha44f, 16'h836c, 16'h8b69, 16'h6a88, 16'h6248, 16'h5a67, 16'h5a67, 16'h5a67, 16'h5a67, 16'h5a68, 16'h6268, 16'h6268, 16'h6288, 16'h72e9, 16'h9c2d, 16'h72e9, 16'h49c5, 16'h1061, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h840, 16'h840, 16'h294, 16'ha44f, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'ha490, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha450, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9ce, 16'h9ce, 16'h9ce, 16'h9ce, 16'h94e, 16'h94e, 16'h94e, 16'h94d, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94d, 16'h94d, 16'h94d, 16'h94d, 16'h94d, 16'h94d, 16'h94e, 16'h93ee, 16'h93ed, 16'h93ee, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93cd, 16'h93cd, 16'h8bcd, 16'h8bcd, 16'h8bcd, 16'h8bac, 16'h5227, 16'h293, 16'h20e2, 16'h20e2, 16'h20e2, 16'h18c1, 16'h840, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h73a, 16'h7b2b, 16'h7b2b, 16'h7b2a, 16'h7b4b, 16'h836c, 16'h838c, 16'h838c, 16'h83ac, 16'h83ac, 16'h8bac, 16'h8bcd, 16'h8bcc, 16'h8bed, 16'h8bed, 16'h94e, 16'h94e, 16'h942e, 16'h942e, 16'h94e, 16'h41c5, 16'h18a1, 16'h212, 16'h3143, 16'h41a5, 16'h4a26, 16'h5a88, 16'h6ba, 16'h734b, 16'h7b8c, 16'h7b8c, 16'h39c6, 16'h1082, 16'h861, 16'h2943, 16'h41e5, 16'h41e5, 16'h41e5, 16'h5226, 16'h3164, 16'h860, 16'h3963, 16'h4184, 16'h3984, 16'h3984, 16'h41a4, 16'h41a4, 16'h3143, 16'h820, 16'h00, 16'h00, 16'h20e3, 16'h3144, 16'h5a47, 16'h5a27, 16'h4a7, 16'h41c6, 16'h3985, 16'h2924, 16'h20e3, 16'h18a2, 16'h861, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h840, 16'h860, 16'h860, 16'h1080, 16'h1081, 16'h1081, 16'h3144, 16'ha490, 16'hb4f1, 16'hacd1, 16'h6ac9, 16'h838, 16'h6aa8, 16'h5a68, 16'h5a67, 16'h5a67, 16'h5a67, 16'h5a67, 16'h6268, 16'h6268, 16'h6268, 16'h6288, 16'h72e9, 16'h9c2e, 16'h739, 16'h49e5, 16'h1061, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h040, 16'h840, 16'h3124, 16'ha44f, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb1, 16'hacb0, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha450, 16'ha450, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha470, 16'ha46f, 16'ha46f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c2e, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9ce, 16'h9ce, 16'h9ce, 16'h9ce, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h93ee, 16'h93ee, 16'h93ee, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ee, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93cd, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93cd, 16'h93cc, 16'h93cd, 16'h93cd, 16'h8b8c, 16'h5227, 16'h293, 16'h20e2, 16'h20e2, 16'h20e2, 16'h18c1, 16'h840, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h732a, 16'h7b4a, 16'h7b4b, 16'h7b4b, 16'h836b, 16'h836c, 16'h838c, 16'h836c, 16'h83ac, 16'h83ac, 16'h83ac, 16'h83ac, 16'h8bcc, 16'h8bcd, 16'h8bed, 16'h8bed, 16'h94e, 16'h94e, 16'h942e, 16'h942e, 16'h7b4b, 16'h732b, 16'h83ac, 16'h8bed, 16'h942e, 16'h9c4f, 16'h942f, 16'h7b4c, 16'h4a27, 16'h3185, 16'h2924, 16'h1081, 16'h841, 16'h040, 16'h861, 16'h1081, 16'h1081, 16'h1081, 16'h1081, 16'h861, 16'h840, 16'h3143, 16'h3984, 16'h3984, 16'h3984, 16'h3984, 16'h3984, 16'h2922, 16'h840, 16'h020, 16'h020, 16'h840, 16'h18a2, 16'h20c2, 16'h1081, 16'h1061, 16'h841, 16'h840, 16'h040, 16'h020, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h860, 16'h860, 16'h860, 16'h1080, 16'h1081, 16'h1081, 16'h1081, 16'h3165, 16'ha490, 16'hb4f1, 16'hacd0, 16'h6288, 16'h7b7, 16'h6aa7, 16'h5a68, 16'h5a67, 16'h5a67, 16'h5a67, 16'h5a67, 16'h6268, 16'h6268, 16'h6268, 16'h6288, 16'h72e9, 16'h9c2d, 16'h739, 16'h41c5, 16'h1061, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h840, 16'h840, 16'h2924, 16'ha44f, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha450, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha46f, 16'ha44f, 16'ha44f, 16'ha46f, 16'ha46f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9ce, 16'h9ce, 16'h9ce, 16'h9ce, 16'h9ce, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94d, 16'h94d, 16'h94d, 16'h93ee, 16'h94e, 16'h93ed, 16'h93ee, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h8bcd, 16'h8b8c, 16'h5227, 16'h293, 16'h212, 16'h20e1, 16'h20e1, 16'h18c1, 16'h840, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h7b2a, 16'h7b2a, 16'h732a, 16'h7b4b, 16'h7b2b, 16'h7b4b, 16'h7b4b, 16'h7b4b, 16'h838c, 16'h838c, 16'h838c, 16'h838c, 16'h838c, 16'h8bcc, 16'h8bcd, 16'h8bed, 16'h94d, 16'h94e, 16'h94e, 16'h942f, 16'h9c2f, 16'h9c4f, 16'h9c4f, 16'h8bad, 16'h7b6c, 16'h6bb, 16'h4a48, 16'h2924, 16'h18a2, 16'h841, 16'h840, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h840, 16'h292, 16'h2923, 16'h213, 16'h20e2, 16'h18c2, 16'h10a1, 16'h1081, 16'h840, 16'h040, 16'h040, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h840, 16'h860, 16'h860, 16'h860, 16'h1080, 16'h1081, 16'h1081, 16'h1081, 16'h3165, 16'ha490, 16'hb4f1, 16'hacd1, 16'h6aa9, 16'h7b7, 16'h6aa7, 16'h5a67, 16'h5a67, 16'h5a67, 16'h5a67, 16'h5a67, 16'h6268, 16'h6267, 16'h6268, 16'h6a88, 16'h72e9, 16'h9c2d, 16'h739, 16'h41e5, 16'h1061, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h040, 16'h840, 16'h2924, 16'h9c6f, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha450, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha46f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4e, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9ce, 16'h94e, 16'h94e, 16'h94e, 16'h9ce, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94d, 16'h94d, 16'h94e, 16'h94d, 16'h93ed, 16'h93ee, 16'h94d, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93cd, 16'h93cd, 16'h93cd, 16'h8bcd, 16'h8bcd, 16'h93cd, 16'h8bcd, 16'h8bcd, 16'h8b8c, 16'h5227, 16'h293, 16'h212, 16'h20e2, 16'h20e2, 16'h18c1, 16'h840, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h7b2a, 16'h6ae9, 16'h73a, 16'h7b4b, 16'h7b2b, 16'h7b4b, 16'h7b4b, 16'h7b4b, 16'h7b4c, 16'h836c, 16'h836c, 16'h836c, 16'h838c, 16'h83ac, 16'h8bcd, 16'h8bed, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h942e, 16'h9c4f, 16'h8bed, 16'h3985, 16'h10a2, 16'h861, 16'h040, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h040, 16'h1081, 16'h840, 16'h840, 16'h860, 16'h860, 16'h840, 16'h040, 16'h040, 16'h020, 16'h020, 16'h020, 16'h020, 16'h040, 16'h020, 16'h020, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h860, 16'h860, 16'h880, 16'h1080, 16'h1081, 16'h1081, 16'h1061, 16'h2924, 16'h9c6f, 16'hb4f1, 16'hacd1, 16'h7b2a, 16'h8327, 16'h6aa7, 16'h5a67, 16'h5a67, 16'h5a67, 16'h5a67, 16'h5a67, 16'h5a68, 16'h6268, 16'h6267, 16'h6a88, 16'h72e9, 16'h9c2d, 16'h739, 16'h49c5, 16'h1061, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h840, 16'h840, 16'h2924, 16'h9c6f, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4e, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9ce, 16'h9ce, 16'h9ce, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94d, 16'h94d, 16'h93ee, 16'h93ee, 16'h93ee, 16'h93ed, 16'h93ed, 16'h93ee, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93cd, 16'h93cd, 16'h8bcd, 16'h8bcd, 16'h8bcd, 16'h8bcd, 16'h8bcd, 16'h8bad, 16'h8b8c, 16'h5227, 16'h293, 16'h212, 16'h211, 16'h20e1, 16'h18c1, 16'h840, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h73a, 16'h6aa8, 16'h739, 16'h732a, 16'h7b2a, 16'h7b2a, 16'h7b4b, 16'h7b4b, 16'h7b4c, 16'h836c, 16'h838c, 16'h83ac, 16'h7b4b, 16'h73b, 16'h7b4b, 16'h8bcd, 16'h94e, 16'h93ee, 16'h8bce, 16'h93ee, 16'h942e, 16'h9c4f, 16'h8bed, 16'h2923, 16'h040, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h861, 16'h2923, 16'h861, 16'h040, 16'h840, 16'h040, 16'h020, 16'h040, 16'h040, 16'h020, 16'h020, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h860, 16'h860, 16'h860, 16'h1080, 16'h1081, 16'h1081, 16'h1061, 16'h18a2, 16'h8bee, 16'hb4d0, 16'hb4d0, 16'h8b8b, 16'h8b48, 16'h6a87, 16'h5a67, 16'h5a67, 16'h5a67, 16'h5a67, 16'h5a67, 16'h5a68, 16'h6268, 16'h6268, 16'h6288, 16'h72e9, 16'h9c2d, 16'h739, 16'h49c5, 16'h1061, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h040, 16'h840, 16'h840, 16'h2924, 16'h9c4f, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb0, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha46f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4e, 16'h9c2e, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9ce, 16'h9ce, 16'h9ce, 16'h94d, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h93ee, 16'h93ee, 16'h93ee, 16'h93ee, 16'h93ed, 16'h93ed, 16'h93ee, 16'h93ee, 16'h93ee, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93cd, 16'h93cd, 16'h93cd, 16'h8bcd, 16'h8bcd, 16'h8bcd, 16'h8bcd, 16'h8bcd, 16'h8bcd, 16'h838c, 16'h5247, 16'h293, 16'h212, 16'h212, 16'h20e2, 16'h18c1, 16'h840, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h73a, 16'h72e9, 16'h7b2a, 16'h7b4b, 16'h7b6b, 16'h7b6b, 16'h836c, 16'h838c, 16'h836c, 16'h838c, 16'h83ac, 16'h83ac, 16'h732b, 16'h6aea, 16'h73a, 16'h838c, 16'h8bed, 16'h8bcd, 16'h8bcd, 16'h93ee, 16'h94e, 16'h942e, 16'h8bed, 16'h2943, 16'h840, 16'h020, 16'h020, 16'h020, 16'h00, 16'h020, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h841, 16'h3144, 16'h1081, 16'h020, 16'h020, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h840, 16'h040, 16'h040, 16'h040, 16'h840, 16'h840, 16'h860, 16'h860, 16'h860, 16'h860, 16'h860, 16'h1061, 16'h7b4c, 16'hb4d1, 16'hacb0, 16'h8bac, 16'h93aa, 16'h6aa7, 16'h5a67, 16'h6267, 16'h6267, 16'h5a68, 16'h5a68, 16'h5a68, 16'h6267, 16'h6267, 16'h6a88, 16'h72e9, 16'h9c2d, 16'h72e9, 16'h49c5, 16'h1061, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h840, 16'h840, 16'h3123, 16'h9c6f, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha46f, 16'ha44f, 16'ha44f, 16'ha46f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9ce, 16'h9ce, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94d, 16'h94e, 16'h94e, 16'h94d, 16'h93ee, 16'h93ee, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93cd, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93cd, 16'h93cd, 16'h8bcd, 16'h8bcd, 16'h8bcd, 16'h8bcd, 16'h8bad, 16'h8bad, 16'h838c, 16'h5227, 16'h213, 16'h20e2, 16'h20e2, 16'h20e2, 16'h18c1, 16'h840, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h73a, 16'h732a, 16'h7b4a, 16'h836b, 16'h836b, 16'h7b4b, 16'h7b4b, 16'h7b6b, 16'h836c, 16'h838c, 16'h83ac, 16'h838c, 16'h732b, 16'h6ae9, 16'h73a, 16'h838c, 16'h8bcd, 16'h8bce, 16'h8bce, 16'h94e, 16'h942f, 16'h9c4f, 16'h94d, 16'h2943, 16'h840, 16'h020, 16'h00, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h841, 16'h3143, 16'h1081, 16'h840, 16'h020, 16'h020, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h840, 16'h840, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h040, 16'h040, 16'h040, 16'h040, 16'h840, 16'h840, 16'h5a89, 16'ha44f, 16'h9c2f, 16'h73a, 16'h9389, 16'h6aa8, 16'h6267, 16'h6267, 16'h6267, 16'h5a68, 16'h5a68, 16'h6268, 16'h6268, 16'h6268, 16'h6a88, 16'h72e9, 16'h9c2d, 16'h739, 16'h49c5, 16'h1061, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h840, 16'h840, 16'h2924, 16'ha46f, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha46f, 16'ha46f, 16'h94e, 16'h7b4b, 16'h838d, 16'h9c4f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9ce, 16'h9ce, 16'h9ce, 16'h94e, 16'h94e, 16'h94e, 16'h94d, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94d, 16'h94d, 16'h94d, 16'h93ed, 16'h93ee, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h8bcd, 16'h8bcd, 16'h8bcd, 16'h8bad, 16'h8bad, 16'h8bad, 16'h8bad, 16'h838c, 16'h5227, 16'h212, 16'h20e2, 16'h20e2, 16'h20e1, 16'h20c1, 16'h840, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h739, 16'h732a, 16'h7b4b, 16'h836b, 16'h7b4b, 16'h732b, 16'h732b, 16'h7b4b, 16'h7b6b, 16'h838c, 16'h838c, 16'h83ad, 16'h7b4b, 16'h73a, 16'h7b4b, 16'h83ac, 16'h8bcd, 16'h93ed, 16'h94e, 16'h942e, 16'h9c4f, 16'h9c4f, 16'h94d, 16'h2943, 16'h840, 16'h00, 16'h020, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h861, 16'h3964, 16'h18a1, 16'h1060, 16'h020, 16'h020, 16'h040, 16'h020, 16'h020, 16'h020, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h040, 16'h040, 16'h840, 16'h860, 16'h41c6, 16'h9c2e, 16'h9c4e, 16'h6267, 16'h7b7, 16'h6aa7, 16'h6267, 16'h6267, 16'h6267, 16'h5a67, 16'h5a68, 16'h6248, 16'h6268, 16'h6268, 16'h6288, 16'h72e9, 16'h9c2d, 16'h739, 16'h41e5, 16'h1061, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h840, 16'h840, 16'h3124, 16'ha44f, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha48f, 16'ha490, 16'ha470, 16'ha470, 16'ha46f, 16'ha46f, 16'h94e, 16'h5228, 16'h3124, 16'h3165, 16'h6289, 16'h9c2e, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9ce, 16'h9ce, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94d, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94d, 16'h93ed, 16'h93ee, 16'h93ee, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h8bcd, 16'h8bcd, 16'h8bcd, 16'h8bad, 16'h8bad, 16'h8bad, 16'h8bad, 16'h838c, 16'h5227, 16'h292, 16'h212, 16'h20e2, 16'h20e1, 16'h18c1, 16'h840, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h73a, 16'h73a, 16'h7b2b, 16'h7b4b, 16'h7b4b, 16'h7b4b, 16'h7b4b, 16'h7b4b, 16'h7b4b, 16'h7b6b, 16'h838c, 16'h83ac, 16'h83ac, 16'h83ac, 16'h8bcd, 16'h8bed, 16'h94d, 16'h94e, 16'h942e, 16'h9c2f, 16'h9c4f, 16'h9c6f, 16'h94e, 16'h3143, 16'h840, 16'h00, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h1061, 16'h4184, 16'h18a1, 16'h1081, 16'h840, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h040, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h840, 16'h840, 16'h840, 16'h840, 16'h3164, 16'ha490, 16'hacb0, 16'h6a88, 16'h7b7, 16'h6a87, 16'h6267, 16'h6267, 16'h6267, 16'h5a68, 16'h5a48, 16'h6268, 16'h6268, 16'h6268, 16'h6288, 16'h72e9, 16'h9c2d, 16'h739, 16'h41e5, 16'h1061, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h840, 16'h840, 16'h3124, 16'ha44f, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacb1, 16'hacb0, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha48f, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha46f, 16'h732b, 16'h3144, 16'h3144, 16'h3124, 16'h3965, 16'h836c, 16'h9c2f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4e, 16'h9c4e, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9ce, 16'h9c2e, 16'h9ce, 16'h9ce, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94d, 16'h94d, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h8bcd, 16'h8bcd, 16'h8bad, 16'h8bac, 16'h8bad, 16'h8bac, 16'h838c, 16'h5227, 16'h293, 16'h20e2, 16'h20e2, 16'h20e1, 16'h18a2, 16'h820, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h739, 16'h73a, 16'h732a, 16'h7b2a, 16'h7b4a, 16'h7b4b, 16'h7b4b, 16'h7b4b, 16'h836b, 16'h838b, 16'h838c, 16'h83ac, 16'h83ac, 16'h8bcd, 16'h8bed, 16'h94e, 16'h942e, 16'h8bed, 16'h94e, 16'h9c2f, 16'h9c4f, 16'h9c6f, 16'h94e, 16'h3143, 16'h840, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h841, 16'h18a2, 16'h41a5, 16'h18a2, 16'h1081, 16'h861, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h040, 16'h040, 16'h040, 16'h020, 16'h040, 16'h040, 16'h040, 16'h040, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h840, 16'h860, 16'h840, 16'h840, 16'h020, 16'h20e3, 16'h9c2e, 16'hacb0, 16'h6288, 16'h837, 16'h6a87, 16'h6247, 16'h6247, 16'h6247, 16'h5a68, 16'h5a67, 16'h6267, 16'h6267, 16'h6268, 16'h6288, 16'h72e9, 16'h9c2d, 16'h739, 16'h49e5, 16'h1061, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h840, 16'h840, 16'h2924, 16'ha44f, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha48f, 16'ha46f, 16'ha46f, 16'ha470, 16'h9c4f, 16'h62a9, 16'h3144, 16'h3144, 16'h3124, 16'h3144, 16'h6269, 16'h8b8d, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c4f, 16'h9c2f, 16'h9c2e, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9ce, 16'h9ce, 16'h9ce, 16'h9ce, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94d, 16'h94d, 16'h94d, 16'h94d, 16'h93ee, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h8bcd, 16'h8bad, 16'h8bad, 16'h8bad, 16'h8bad, 16'h838c, 16'h5227, 16'h213, 16'h212, 16'h20e2, 16'h20e2, 16'h18a2, 16'h840, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h739, 16'h7329, 16'h7b2a, 16'h7b2a, 16'h7b2a, 16'h7b4b, 16'h7b6b, 16'h836b, 16'h832b, 16'h836b, 16'h83ac, 16'h8bcc, 16'h8bcd, 16'h93cd, 16'h93ed, 16'h9bac, 16'h9c2e, 16'h7b4b, 16'h83ac, 16'h9c2f, 16'h9c4f, 16'h9c6f, 16'h94e, 16'h3143, 16'h840, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h861, 16'h2923, 16'h3143, 16'h49c5, 16'h20c2, 16'h10a1, 16'h1081, 16'h020, 16'h020, 16'h840, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h040, 16'h040, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h840, 16'h860, 16'h861, 16'h860, 16'h820, 16'h020, 16'h020, 16'h1082, 16'h8bcd, 16'hacb0, 16'h6288, 16'h838, 16'h6a88, 16'h6248, 16'h5a48, 16'h6248, 16'h5a47, 16'h5a67, 16'h5a67, 16'h6267, 16'h6267, 16'h6288, 16'h72e9, 16'h9c2e, 16'h739, 16'h49c5, 16'h1061, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h840, 16'h840, 16'h3124, 16'ha44f, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha46f, 16'h9c4f, 16'h5248, 16'h3964, 16'h3144, 16'h2923, 16'h3964, 16'h527, 16'h834c, 16'h9c2e, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9ce, 16'h9ce, 16'h9ce, 16'h9ce, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94d, 16'h94e, 16'h94d, 16'h94d, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h8bcd, 16'h93cd, 16'h93cd, 16'h8bcc, 16'h8bac, 16'h8bad, 16'h8bad, 16'h8bad, 16'h836c, 16'h5227, 16'h292, 16'h212, 16'h20e1, 16'h20e2, 16'h18c1, 16'h840, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h739, 16'h7b2a, 16'h7b2a, 16'h7aea, 16'h72c9, 16'h7b2b, 16'h7b4b, 16'h834b, 16'h7ac9, 16'h7b2a, 16'h838c, 16'h83ac, 16'h8bcc, 16'h93ac, 16'h8a89, 16'h8a7, 16'h9bcd, 16'h73a, 16'h7b6b, 16'h9c4f, 16'h9c4f, 16'h9c6f, 16'h94e, 16'h3143, 16'h840, 16'h020, 16'h020, 16'h020, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h820, 16'h1061, 16'h1882, 16'h49a5, 16'h20c2, 16'h18a1, 16'h1081, 16'h840, 16'h020, 16'h840, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h840, 16'h840, 16'h840, 16'h18c2, 16'h18c1, 16'h840, 16'h020, 16'h020, 16'h841, 16'h7b4c, 16'hacb0, 16'h6268, 16'h838, 16'h6a88, 16'h6247, 16'h5a47, 16'h6247, 16'h5a47, 16'h5a67, 16'h5a67, 16'h5a67, 16'h6267, 16'h6288, 16'h72e9, 16'h9cd, 16'h739, 16'h49e5, 16'h1061, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h840, 16'h840, 16'h314, 16'ha44f, 16'hb4d1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'h9c2f, 16'h5a48, 16'h3984, 16'h3143, 16'h213, 16'h3964, 16'h4165, 16'h6249, 16'h8bad, 16'h9c4e, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9ce, 16'h94e, 16'h94e, 16'h94e, 16'h94d, 16'h94d, 16'h94e, 16'h94e, 16'h94d, 16'h93ee, 16'h93ee, 16'h93ed, 16'h94d, 16'h94d, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h8bcd, 16'h8bcd, 16'h8bcd, 16'h8bcd, 16'h8bcd, 16'h8bcd, 16'h8bad, 16'h8bad, 16'h8bad, 16'h8bad, 16'h8bad, 16'h836c, 16'h5227, 16'h293, 16'h20e2, 16'h20e2, 16'h20e2, 16'h18c1, 16'h840, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h72e9, 16'h7b2a, 16'h7b2a, 16'h7ac9, 16'h7ac9, 16'h7b4b, 16'h7b4b, 16'h7b4b, 16'h7ac9, 16'h832a, 16'h8bac, 16'h83ac, 16'h8bcc, 16'h93cc, 16'h8a47, 16'h89e7, 16'h9bcd, 16'h732a, 16'h7b6b, 16'h942f, 16'h9c4f, 16'h9c6f, 16'h94e, 16'h3143, 16'h840, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h841, 16'h49a5, 16'h20c2, 16'h18a1, 16'h18a1, 16'h840, 16'h00, 16'h840, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h040, 16'h880, 16'h860, 16'h040, 16'h020, 16'h840, 16'h212, 16'h18e1, 16'h840, 16'h020, 16'h020, 16'h821, 16'h6aea, 16'hacb0, 16'h5a67, 16'h7b7, 16'h6a87, 16'h5a47, 16'h5a47, 16'h6247, 16'h5a47, 16'h5a67, 16'h5a47, 16'h6267, 16'h6267, 16'h6287, 16'h72e9, 16'h9ce, 16'h73a, 16'h41e5, 16'h1061, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h840, 16'h3123, 16'h9c4f, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb0, 16'hacb0, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb1, 16'hacb1, 16'hacb0, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha48f, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha46f, 16'ha46f, 16'h9c2f, 16'h5a68, 16'h3964, 16'h2923, 16'h18c2, 16'h20e2, 16'h2924, 16'h3965, 16'h62a9, 16'h9c2e, 16'h9c2f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9ce, 16'h9c2e, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94d, 16'h94e, 16'h93ee, 16'h93ee, 16'h93ed, 16'h93ed, 16'h94d, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h8bcd, 16'h8bcd, 16'h8bad, 16'h8bcd, 16'h8bcd, 16'h8bcd, 16'h8bcd, 16'h8bad, 16'h8bad, 16'h8bac, 16'h8bad, 16'h8b8d, 16'h836c, 16'h5227, 16'h213, 16'h20e2, 16'h20e2, 16'h20c2, 16'h18a1, 16'h820, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h72e9, 16'h7b2a, 16'h7b2a, 16'h7ac9, 16'h7ae9, 16'h834b, 16'h7b4a, 16'h7b4b, 16'h82a9, 16'h832b, 16'h836c, 16'h838c, 16'h8bac, 16'h93cc, 16'h8a67, 16'h927, 16'h9bcd, 16'h7b4b, 16'h7b4b, 16'h942f, 16'h9c4f, 16'h9c4f, 16'h94e, 16'h3143, 16'h840, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h821, 16'h49a5, 16'h28e2, 16'h18a2, 16'h18a2, 16'h861, 16'h00, 16'h841, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h00, 16'h020, 16'h840, 16'h840, 16'h18e2, 16'h18c1, 16'h840, 16'h020, 16'h020, 16'h020, 16'h5a69, 16'hacb0, 16'h5a67, 16'h838, 16'h6a87, 16'h5a47, 16'h5a47, 16'h6247, 16'h5a67, 16'h5a47, 16'h5a47, 16'h6267, 16'h6268, 16'h6288, 16'h72e9, 16'h9c2e, 16'h73a, 16'h41e5, 16'h1061, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h840, 16'h2923, 16'h9c4f, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'h9c4f, 16'h6aaa, 16'h3965, 16'h3124, 16'h18a2, 16'h10a2, 16'h18c2, 16'h213, 16'h39a5, 16'h8bcd, 16'h9c2f, 16'h9c4f, 16'h9c2e, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h94e, 16'h9ce, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94d, 16'h93ed, 16'h93ee, 16'h93ee, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h8bcd, 16'h8bcd, 16'h8bcd, 16'h8bad, 16'h8bad, 16'h8bad, 16'h8bad, 16'h8bad, 16'h8bad, 16'h8bad, 16'h8bad, 16'h8bac, 16'h8bac, 16'h8b8d, 16'h836c, 16'h5227, 16'h213, 16'h20e2, 16'h20e2, 16'h20e2, 16'h18c1, 16'h840, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h7ba, 16'h7b2a, 16'h7b2a, 16'h7ac9, 16'h7ae9, 16'h834b, 16'h7b4b, 16'h7b2a, 16'h7aa9, 16'h834b, 16'h838c, 16'h838c, 16'h8bac, 16'h93cc, 16'h8a47, 16'h91a6, 16'ha3ad, 16'h836b, 16'h7b4b, 16'h942e, 16'h9c4f, 16'h9c4f, 16'h8cd, 16'h3163, 16'h840, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h821, 16'h49a5, 16'h293, 16'h20c2, 16'h20a2, 16'h1061, 16'h00, 16'h841, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h00, 16'h00, 16'h00, 16'h020, 16'h840, 16'h840, 16'h10a1, 16'h1081, 16'h820, 16'h020, 16'h020, 16'h00, 16'h4a7, 16'ha490, 16'h5a47, 16'h837, 16'h6a88, 16'h5a47, 16'h5a47, 16'h5a47, 16'h5a47, 16'h5a47, 16'h5a47, 16'h6267, 16'h6268, 16'h6288, 16'h72e9, 16'h9c2e, 16'h73a, 16'h41e5, 16'h1061, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h840, 16'h3124, 16'h9c4f, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha470, 16'h9c4f, 16'h732b, 16'h3984, 16'h3964, 16'h20e2, 16'h1881, 16'h18a2, 16'h293, 16'h294, 16'h7b4b, 16'h9c2e, 16'h9c4e, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9ce, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94d, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94d, 16'h94d, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h8bcd, 16'h8bcd, 16'h8bcd, 16'h8bcd, 16'h8bcc, 16'h8bcc, 16'h8bcc, 16'h8bad, 16'h8bad, 16'h8bad, 16'h8bad, 16'h8bac, 16'h8bac, 16'h8bac, 16'h8bac, 16'h8bac, 16'h8b8d, 16'h836c, 16'h5227, 16'h293, 16'h20e2, 16'h20e2, 16'h20e2, 16'h18c1, 16'h840, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h7ba, 16'h7b2a, 16'h7b2a, 16'h7aa9, 16'h7ba, 16'h834b, 16'h7b4b, 16'h7b4a, 16'h82a9, 16'h834b, 16'h838c, 16'h838c, 16'h8bac, 16'h93ad, 16'h8a47, 16'h8965, 16'ha3ad, 16'h83ac, 16'h7b6b, 16'h942e, 16'h9c4f, 16'h9c4f, 16'h94d, 16'h3163, 16'h840, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h820, 16'h49c5, 16'h2923, 16'h20e2, 16'h18c2, 16'h1061, 16'h00, 16'h841, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h00, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h00, 16'h00, 16'h00, 16'h3985, 16'ha46f, 16'h5a47, 16'h7ae7, 16'h6a87, 16'h5a67, 16'h5a67, 16'h6247, 16'h5a47, 16'h5a47, 16'h5a47, 16'h5a48, 16'h6267, 16'h6288, 16'h72e9, 16'h9c2e, 16'h7b2a, 16'h41e5, 16'h1061, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h840, 16'h2924, 16'h9c4f, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha44f, 16'h8bad, 16'h41a5, 16'h41a4, 16'h3143, 16'h18a2, 16'h18a2, 16'h213, 16'h20e3, 16'h6ac9, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9ce, 16'h9ce, 16'h9ce, 16'h9ce, 16'h9ce, 16'h9ce, 16'h9ce, 16'h94e, 16'h94d, 16'h94d, 16'h94e, 16'h94d, 16'h94d, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93cd, 16'h93ed, 16'h93ed, 16'h93cd, 16'h8bcd, 16'h93cd, 16'h93cd, 16'h8bcd, 16'h8bcd, 16'h8bcc, 16'h8bcc, 16'h8bac, 16'h8bad, 16'h8bad, 16'h8bad, 16'h8bad, 16'h8bac, 16'h8bac, 16'h8bac, 16'h8bac, 16'h8b8d, 16'h836c, 16'h526, 16'h212, 16'h20e2, 16'h20e2, 16'h20e2, 16'h18c1, 16'h840, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h7ba, 16'h7b2a, 16'h7b2a, 16'h7aa9, 16'h7aea, 16'h7b2b, 16'h834b, 16'h834a, 16'h82a9, 16'h834b, 16'h8b8c, 16'h838c, 16'h838c, 16'h8bac, 16'h8a27, 16'h8965, 16'h9b4c, 16'h8bcc, 16'h838b, 16'h942e, 16'h9c4f, 16'h9c4f, 16'h8cd, 16'h3163, 16'h840, 16'h020, 16'h020, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h820, 16'h49c5, 16'h3123, 16'h20e2, 16'h18c2, 16'h1081, 16'h00, 16'h861, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h00, 16'h00, 16'h820, 16'h841, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h3144, 16'h9c4e, 16'h5227, 16'h7ac7, 16'h6a88, 16'h5a47, 16'h6247, 16'h6247, 16'h5a47, 16'h5a47, 16'h5a47, 16'h6268, 16'h6268, 16'h6288, 16'h72e9, 16'h9c2e, 16'h732a, 16'h41c5, 16'h1061, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h840, 16'h2923, 16'ha44f, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha44f, 16'h94e, 16'h527, 16'h4184, 16'h41a4, 16'h20e2, 16'h18a2, 16'h20c2, 16'h20c3, 16'h5a48, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9ce, 16'h9ce, 16'h9ce, 16'h9ce, 16'h9ce, 16'h94e, 16'h94e, 16'h94e, 16'h94d, 16'h94d, 16'h94d, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h8bcd, 16'h8bcd, 16'h8bcc, 16'h8bcc, 16'h8bcc, 16'h8bcc, 16'h8bad, 16'h8bad, 16'h8bac, 16'h8bac, 16'h8bad, 16'h8bac, 16'h8bac, 16'h8bac, 16'h8bac, 16'h8b8c, 16'h836b, 16'h526, 16'h292, 16'h20e2, 16'h20e2, 16'h20c2, 16'h18a1, 16'h840, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h7b2a, 16'h7b4a, 16'h7b2a, 16'h7aa9, 16'h7ba, 16'h7b4b, 16'h7b4b, 16'h832a, 16'h7aa9, 16'h832b, 16'h838c, 16'h838c, 16'h838c, 16'h8b8c, 16'h8a47, 16'h8964, 16'h93b, 16'h8bcd, 16'h83ac, 16'h942e, 16'h9c4f, 16'h9c4f, 16'h94e, 16'h3163, 16'h040, 16'h020, 16'h020, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h841, 16'h49c5, 16'h3124, 16'h20e3, 16'h20c3, 16'h1081, 16'h00, 16'h861, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h841, 16'h213, 16'h3144, 16'h18c2, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h20e3, 16'h9c2e, 16'h5a27, 16'h7aa7, 16'h6a88, 16'h5a47, 16'h6247, 16'h5a47, 16'h5a48, 16'h5a47, 16'h5a48, 16'h6268, 16'h6268, 16'h6288, 16'h72c9, 16'h9c2e, 16'h7b2a, 16'h41c5, 16'h1061, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h840, 16'h2923, 16'ha44f, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha470, 16'ha46f, 16'ha470, 16'ha46f, 16'ha44f, 16'h9c4f, 16'h6ac9, 16'h3964, 16'h41a4, 16'h2923, 16'h18a2, 16'h20c2, 16'h18c2, 16'h4a7, 16'h94e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9ce, 16'h9ce, 16'h9ce, 16'h9ce, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94d, 16'h94d, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h8bcd, 16'h8bcd, 16'h8bcd, 16'h8bad, 16'h8bcc, 16'h8bad, 16'h8bad, 16'h8bad, 16'h8bac, 16'h8bac, 16'h8bac, 16'h8bac, 16'h8bac, 16'h8bac, 16'h8bac, 16'h8bac, 16'h8b8c, 16'h834c, 16'h526, 16'h293, 16'h20e2, 16'h20e2, 16'h20c2, 16'h18a1, 16'h820, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h72ea, 16'h7b2a, 16'h7b2a, 16'h7a88, 16'h7ba, 16'h834b, 16'h834b, 16'h834b, 16'h7aa9, 16'h7ba, 16'h838c, 16'h836c, 16'h838c, 16'h8b8b, 16'h8227, 16'h8964, 16'h92ea, 16'h93ed, 16'h8bcc, 16'h942e, 16'h9c4f, 16'h9c4f, 16'h94d, 16'h3163, 16'h840, 16'h020, 16'h020, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h1081, 16'h51e6, 16'h3144, 16'h20e3, 16'h20e3, 16'h1081, 16'h00, 16'h861, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h040, 16'h040, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h841, 16'h3164, 16'h3984, 16'h20e2, 16'h820, 16'h00, 16'h00, 16'h00, 16'h020, 16'h840, 16'h820, 16'h020, 16'h18c2, 16'h94e, 16'h5a47, 16'h72a6, 16'h6a87, 16'h5a47, 16'h5a47, 16'h5a47, 16'h5a48, 16'h5a47, 16'h5a47, 16'h5a67, 16'h6268, 16'h6a88, 16'h72c9, 16'h9c2e, 16'h7b4a, 16'h49e5, 16'h1061, 16'h00, 16'h821, 16'h820, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h840, 16'h2923, 16'ha44f, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha48f, 16'ha46f, 16'ha470, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha44f, 16'ha44f, 16'h8bad, 16'h41a5, 16'h3144, 16'h20e3, 16'h18a2, 16'h18c2, 16'h18c2, 16'h4a7, 16'h94e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9ce, 16'h9ce, 16'h94e, 16'h94e, 16'h94d, 16'h94e, 16'h94e, 16'h94d, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93cd, 16'h93ed, 16'h93cd, 16'h93cd, 16'h93cd, 16'h8bcd, 16'h8bcd, 16'h8bcc, 16'h8bcc, 16'h8bcd, 16'h8bad, 16'h8bac, 16'h8bac, 16'h8bad, 16'h8bac, 16'h8bac, 16'h8bac, 16'h8bac, 16'h8bac, 16'h8bac, 16'h8bac, 16'h8bac, 16'h8b8c, 16'h8b8c, 16'h836b, 16'h526, 16'h292, 16'h212, 16'h20e1, 16'h20e1, 16'h18c1, 16'h840, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h7b2a, 16'h7b2b, 16'h7b2a, 16'h7a89, 16'h7ba, 16'h7b4b, 16'h7b4b, 16'h7b2b, 16'h7aa9, 16'h7ba, 16'h838c, 16'h838c, 16'h838c, 16'h8b8c, 16'h82a8, 16'h8a27, 16'h932b, 16'h93ed, 16'h94d, 16'h942e, 16'h9c4f, 16'h9c4f, 16'h94e, 16'h3183, 16'h840, 16'h020, 16'h020, 16'h020, 16'h00, 16'h020, 16'h00, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h1061, 16'h49c5, 16'h3144, 16'h213, 16'h20e3, 16'h10a2, 16'h020, 16'h861, 16'h840, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h040, 16'h040, 16'h040, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h840, 16'h2943, 16'h3164, 16'h212, 16'h820, 16'h00, 16'h00, 16'h00, 16'h840, 16'h10a1, 16'h18c2, 16'h18c2, 16'h18c2, 16'h7b4b, 16'h5227, 16'h72a6, 16'h6a87, 16'h5a47, 16'h5a47, 16'h5a47, 16'h5a47, 16'h5a47, 16'h5a48, 16'h5a48, 16'h6268, 16'h6288, 16'h72c9, 16'h9c2e, 16'h7b4b, 16'h41e5, 16'h1061, 16'h00, 16'h020, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h840, 16'h3123, 16'ha44f, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'hac90, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha46f, 16'ha470, 16'ha470, 16'ha44f, 16'ha44f, 16'ha46f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c2f, 16'h62a9, 16'h293, 16'h18c3, 16'h18a2, 16'h18c2, 16'h18c2, 16'h5227, 16'h9ce, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9ce, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94d, 16'h94d, 16'h94e, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ec, 16'h93ec, 16'h93cd, 16'h8bed, 16'h93cd, 16'h8bcd, 16'h8bcd, 16'h8bcd, 16'h8bcd, 16'h8bcd, 16'h8bad, 16'h8bac, 16'h8bac, 16'h8bac, 16'h8bac, 16'h8bac, 16'h8bac, 16'h8bac, 16'h8bac, 16'h8b8c, 16'h8b8c, 16'h8bac, 16'h8bac, 16'h8b8c, 16'h834b, 16'h4a6, 16'h28e3, 16'h20e2, 16'h20e2, 16'h20e1, 16'h18c2, 16'h820, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h73a, 16'h73b, 16'h7ba, 16'h7aa8, 16'h7ae9, 16'h7b2a, 16'h732b, 16'h7b2b, 16'h7ac9, 16'h7b2a, 16'h7b6b, 16'h838c, 16'h838b, 16'h8bac, 16'h8bac, 16'h8bcd, 16'h93ed, 16'h94e, 16'h94e, 16'h942e, 16'h942f, 16'h9c2f, 16'h8bed, 16'h3163, 16'h840, 16'h020, 16'h020, 16'h020, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h820, 16'h4185, 16'h3964, 16'h213, 16'h20e3, 16'h18a2, 16'h020, 16'h861, 16'h840, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h040, 16'h040, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h840, 16'h212, 16'h212, 16'h18c2, 16'h841, 16'h00, 16'h00, 16'h00, 16'h00, 16'h820, 16'h861, 16'h1061, 16'h841, 16'h18c3, 16'h20a2, 16'h72a6, 16'h6a87, 16'h5a47, 16'h5a47, 16'h5a47, 16'h5a47, 16'h5a47, 16'h5a47, 16'h6248, 16'h6268, 16'h6a68, 16'h72c9, 16'h9c4e, 16'h836b, 16'h49e5, 16'h1061, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h840, 16'h3124, 16'h9c4f, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'hac90, 16'hac90, 16'hac90, 16'ha48f, 16'ha470, 16'ha470, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h8bcd, 16'h49e6, 16'h213, 16'h20e3, 16'h20e3, 16'h213, 16'h62c9, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9ce, 16'h9c2e, 16'h9ce, 16'h9ce, 16'h9ce, 16'h94e, 16'h94e, 16'h94d, 16'h94d, 16'h94d, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h8bcd, 16'h8bcd, 16'h8bcd, 16'h8bcd, 16'h8bcd, 16'h8bcc, 16'h8bcc, 16'h8bad, 16'h8bad, 16'h8bac, 16'h8bac, 16'h8bac, 16'h8bac, 16'h8bac, 16'h8bac, 16'h8bac, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h834b, 16'h526, 16'h212, 16'h20e2, 16'h20e1, 16'h20e1, 16'h18c2, 16'h840, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h73a, 16'h73a, 16'h7ba, 16'h7ae9, 16'h7b2a, 16'h7b4b, 16'h7b4b, 16'h7b6b, 16'h836b, 16'h838c, 16'h838c, 16'h838c, 16'h83ac, 16'h8bad, 16'h8bcd, 16'h8bed, 16'h93ed, 16'h94e, 16'h94e, 16'h942e, 16'h942f, 16'h9c2f, 16'h8cd, 16'h3164, 16'h840, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h00, 16'h00, 16'h020, 16'h4184, 16'h3984, 16'h2923, 16'h213, 16'h18a2, 16'h020, 16'h861, 16'h840, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h040, 16'h040, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h841, 16'h020, 16'h00, 16'h00, 16'h00, 16'h020, 16'h020, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h040, 16'h1061, 16'h6a85, 16'h6a87, 16'h5a47, 16'h5a47, 16'h5a47, 16'h5a47, 16'h5a47, 16'h5a47, 16'h6248, 16'h6268, 16'h6a88, 16'h72c9, 16'h9c4e, 16'h836b, 16'h49e5, 16'h1061, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h840, 16'h2924, 16'h9c4f, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'hac90, 16'hac90, 16'hac90, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4e, 16'h7b4b, 16'h41c5, 16'h293, 16'h293, 16'h41c6, 16'h838c, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9ce, 16'h9ce, 16'h9ce, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94d, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93cd, 16'h93cd, 16'h93ed, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h8bcd, 16'h8bcd, 16'h8bcd, 16'h8bcd, 16'h8bcd, 16'h8bad, 16'h8bad, 16'h8bad, 16'h8bad, 16'h8bac, 16'h8bac, 16'h8bac, 16'h8b8c, 16'h8bac, 16'h8bac, 16'h8bac, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h838c, 16'h836c, 16'h834b, 16'h4a6, 16'h212, 16'h20e2, 16'h20e1, 16'h20e1, 16'h18c1, 16'h820, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h7b2b, 16'h7b4a, 16'h7b4b, 16'h7b4b, 16'h7b6b, 16'h7b6b, 16'h7b6b, 16'h838b, 16'h838b, 16'h838c, 16'h838c, 16'h838c, 16'h83ac, 16'h83ac, 16'h8bcd, 16'h8bcd, 16'h8bed, 16'h93ee, 16'h94e, 16'h94e, 16'h942e, 16'h9c2e, 16'h8bed, 16'h3184, 16'h840, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h3964, 16'h3964, 16'h2923, 16'h213, 16'h18c2, 16'h020, 16'h861, 16'h840, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h040, 16'h040, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h840, 16'h6a86, 16'h6a87, 16'h5a47, 16'h5a47, 16'h5a47, 16'h5a47, 16'h5a47, 16'h5a47, 16'h5a48, 16'h6248, 16'h6288, 16'h72c9, 16'h9c2e, 16'h836b, 16'h49e5, 16'h1061, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h840, 16'h2924, 16'h9c4f, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'hac90, 16'hac90, 16'hac90, 16'ha490, 16'ha470, 16'ha46f, 16'ha470, 16'ha470, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4e, 16'h9c4e, 16'h838b, 16'h5a67, 16'h526, 16'h73a, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9ce, 16'h9ce, 16'h9ce, 16'h9ce, 16'h9ce, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h93ee, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h8bcd, 16'h8bcd, 16'h8bcd, 16'h8bcd, 16'h8bac, 16'h8bad, 16'h8bad, 16'h8bad, 16'h8bad, 16'h8bac, 16'h8bac, 16'h8bac, 16'h8b8c, 16'h8bac, 16'h8b8c, 16'h8b8c, 16'h838c, 16'h838c, 16'h8b8c, 16'h838c, 16'h838c, 16'h834b, 16'h4a6, 16'h212, 16'h20e2, 16'h20e2, 16'h20e1, 16'h18a1, 16'h820, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h7b4b, 16'h7b4b, 16'h7b4b, 16'h7b4b, 16'h7b6b, 16'h7b6b, 16'h7b6b, 16'h836b, 16'h838c, 16'h838c, 16'h838c, 16'h838c, 16'h838c, 16'h83ac, 16'h8bcc, 16'h8bec, 16'h8bed, 16'h94d, 16'h94e, 16'h94e, 16'h942e, 16'h9c2e, 16'h8bed, 16'h3184, 16'h840, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h040, 16'h840, 16'h840, 16'h840, 16'h840, 16'h860, 16'h1081, 16'h41a4, 16'h3984, 16'h293, 16'h293, 16'h18c2, 16'h020, 16'h861, 16'h840, 16'h020, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h840, 16'h841, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h840, 16'h6a66, 16'h6a87, 16'h5a47, 16'h5a47, 16'h5a47, 16'h5a47, 16'h5a47, 16'h5a47, 16'h5a47, 16'h5a67, 16'h6268, 16'h72c9, 16'h9c2e, 16'h836b, 16'h49c5, 16'h1061, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h840, 16'h2924, 16'h9c4f, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'hac90, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha44f, 16'ha46f, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h94e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9ce, 16'h9ce, 16'h9ce, 16'h9ce, 16'h9ce, 16'h94d, 16'h94e, 16'h93ee, 16'h94d, 16'h94d, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93ed, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h8bcd, 16'h8bcd, 16'h8bad, 16'h8bad, 16'h8bad, 16'h8bad, 16'h8bad, 16'h8bad, 16'h8bad, 16'h8bac, 16'h8bac, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h838c, 16'h838c, 16'h7b4b, 16'h49e6, 16'h292, 16'h20e2, 16'h20e2, 16'h20e1, 16'h18a1, 16'h820, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h7b2b, 16'h7b4b, 16'h7b4b, 16'h7b4b, 16'h7b4c, 16'h7b4c, 16'h7b6b, 16'h836b, 16'h836c, 16'h838c, 16'h838c, 16'h838c, 16'h838c, 16'h83ad, 16'h8bcd, 16'h8bcd, 16'h8bed, 16'h94d, 16'h94d, 16'h94e, 16'h942e, 16'h942e, 16'h8bed, 16'h3984, 16'h840, 16'h020, 16'h040, 16'h840, 16'h860, 16'h860, 16'h1080, 16'h18c1, 16'h212, 16'h3143, 16'h39a4, 16'h4a5, 16'h5a87, 16'h72e8, 16'h6aa7, 16'h4184, 16'h2923, 16'h2923, 16'h18e2, 16'h020, 16'h861, 16'h841, 16'h020, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h840, 16'h10a2, 16'h840, 16'h020, 16'h020, 16'h020, 16'h020, 16'h840, 16'h6a66, 16'h6a87, 16'h5a47, 16'h5a47, 16'h5a47, 16'h5a47, 16'h5a47, 16'h5a47, 16'h5a47, 16'h5a67, 16'h6268, 16'h72c9, 16'h9c2e, 16'h836b, 16'h49c5, 16'h1061, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h020, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h840, 16'h2924, 16'ha46f, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha46f, 16'ha470, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9ce, 16'h9ce, 16'h9ce, 16'h9ce, 16'h9cd, 16'h94d, 16'h94d, 16'h93ed, 16'h93ed, 16'h94d, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93cd, 16'h93ed, 16'h93ed, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h8bcd, 16'h8bcd, 16'h8bad, 16'h8bad, 16'h8bad, 16'h8bad, 16'h8bad, 16'h8bad, 16'h8bac, 16'h8bac, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h836c, 16'h836c, 16'h834b, 16'h49e6, 16'h292, 16'h20e1, 16'h20e2, 16'h20e1, 16'h18a2, 16'h820, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h7b4a, 16'h7b4b, 16'h7b4a, 16'h7b4b, 16'h7b4b, 16'h7b6b, 16'h836b, 16'h836b, 16'h836c, 16'h836c, 16'h838c, 16'h838c, 16'h83ac, 16'h83ac, 16'h8bad, 16'h8bcd, 16'h8bed, 16'h8bed, 16'h94e, 16'h94e, 16'h942e, 16'h942e, 16'h8bed, 16'h3984, 16'h10a1, 16'h18e1, 16'h2922, 16'h3984, 16'h4a5, 16'h5a87, 16'h6ae9, 16'h7b6b, 16'h83ac, 16'h93ed, 16'h942d, 16'h9c2d, 16'h9c2c, 16'h94c, 16'h7ae8, 16'h4184, 16'h2923, 16'h2923, 16'h18e2, 16'h020, 16'h861, 16'h841, 16'h020, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h841, 16'h1082, 16'h840, 16'h020, 16'h020, 16'h020, 16'h020, 16'h840, 16'h6a45, 16'h6a87, 16'h5a47, 16'h5a47, 16'h5a47, 16'h5a47, 16'h5a47, 16'h5a47, 16'h5a47, 16'h6247, 16'h6268, 16'h6ac9, 16'h9cd, 16'h7b6b, 16'h41c5, 16'h1061, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h040, 16'h840, 16'h3124, 16'ha44f, 16'hb4d1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha470, 16'ha490, 16'ha490, 16'ha470, 16'ha46f, 16'ha450, 16'ha46f, 16'ha46f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9ce, 16'h9ce, 16'h9ce, 16'h9cd, 16'h94d, 16'h94d, 16'h93ed, 16'h94d, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93cd, 16'h93cd, 16'h93ed, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h8bcd, 16'h8bcd, 16'h8bcd, 16'h8bad, 16'h8bad, 16'h8bad, 16'h8bad, 16'h8bad, 16'h8bad, 16'h8bad, 16'h8bac, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h838c, 16'h8b8c, 16'h838c, 16'h8b6c, 16'h834b, 16'h49e6, 16'h212, 16'h20e1, 16'h20e2, 16'h20e1, 16'h18a1, 16'h820, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h7b2b, 16'h7b4b, 16'h7b4b, 16'h7b4b, 16'h7b4b, 16'h7b6b, 16'h836b, 16'h836b, 16'h836b, 16'h836c, 16'h838c, 16'h838c, 16'h838c, 16'h83ac, 16'h83ac, 16'h8bcc, 16'h8bed, 16'h8bed, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h732a, 16'h732a, 16'h83ab, 16'h8bec, 16'h942e, 16'h9c4e, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4e, 16'h9c2d, 16'h9c2d, 16'h9c2d, 16'h7b9, 16'h41a5, 16'h2924, 16'h2924, 16'h18e2, 16'h020, 16'h861, 16'h841, 16'h020, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h840, 16'h820, 16'h020, 16'h020, 16'h020, 16'h020, 16'h861, 16'h1061, 16'h6a65, 16'h6a87, 16'h5a47, 16'h5a47, 16'h5a47, 16'h5a47, 16'h5a47, 16'h5a47, 16'h5a47, 16'h5a47, 16'h6267, 16'h6ac9, 16'h9cd, 16'h7b4b, 16'h41e5, 16'h1081, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h040, 16'h840, 16'h3124, 16'ha44f, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha450, 16'ha46f, 16'ha46f, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9ce, 16'h9ce, 16'h9ce, 16'h9ce, 16'h9cd, 16'h94d, 16'h93ee, 16'h94d, 16'h94d, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h8bcd, 16'h8bcd, 16'h8bcd, 16'h8bcd, 16'h8bcc, 16'h8bad, 16'h8bad, 16'h8bad, 16'h8bac, 16'h8bac, 16'h8bad, 16'h8bac, 16'h8bac, 16'h8b8d, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8b, 16'h8b8b, 16'h8b8b, 16'h838c, 16'h8b6c, 16'h7b4b, 16'h4a6, 16'h212, 16'h20e2, 16'h20e2, 16'h20e1, 16'h18a1, 16'h820, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h7b2b, 16'h7b4b, 16'h7b4b, 16'h7b4b, 16'h7b4b, 16'h7b6a, 16'h7b6b, 16'h836b, 16'h836b, 16'h838b, 16'h838c, 16'h838c, 16'h836c, 16'h7b4b, 16'h7b4b, 16'h838c, 16'h8bcd, 16'h8bed, 16'h8bee, 16'h8bee, 16'h8bcd, 16'h94e, 16'h94e, 16'h942e, 16'h942e, 16'h9c4e, 16'h9c4e, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4e, 16'h9c2d, 16'h9c2d, 16'h9c4e, 16'h9c2e, 16'h7ba, 16'h41a4, 16'h3143, 16'h2924, 16'h20e3, 16'h020, 16'h861, 16'h861, 16'h020, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h820, 16'h00, 16'h00, 16'h00, 16'h00, 16'h820, 16'h39a5, 16'h3964, 16'h6a66, 16'h6a67, 16'h5a47, 16'h5a47, 16'h5a47, 16'h5a47, 16'h5a47, 16'h5a47, 16'h5a47, 16'h5a47, 16'h6268, 16'h6ac9, 16'h9cd, 16'h7b4b, 16'h41c5, 16'h1081, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h840, 16'h3124, 16'ha46f, 16'hacd1, 16'hacd1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha470, 16'ha46f, 16'ha470, 16'ha470, 16'ha46f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9ce, 16'h9ce, 16'h9ce, 16'h9ce, 16'h9cd, 16'h94d, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cc, 16'h93cd, 16'h8bcd, 16'h8bcd, 16'h8bcd, 16'h8bad, 16'h8bcd, 16'h8bac, 16'h8bac, 16'h8bad, 16'h8bac, 16'h8bac, 16'h8bac, 16'h8bad, 16'h8bac, 16'h8bac, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8b, 16'h838b, 16'h8b6c, 16'h836c, 16'h8b6b, 16'h7b4b, 16'h4a6, 16'h212, 16'h20e2, 16'h20c2, 16'h20e1, 16'h18a1, 16'h820, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h7b2a, 16'h7b2b, 16'h7b4b, 16'h7b4b, 16'h7b6b, 16'h836b, 16'h836b, 16'h7b6b, 16'h836c, 16'h838c, 16'h838c, 16'h838c, 16'h73a, 16'h62a9, 16'h62a9, 16'h732b, 16'h83ac, 16'h8bcd, 16'h8bad, 16'h8bad, 16'h8bac, 16'h93ed, 16'h93ee, 16'h942e, 16'h9c2e, 16'h9c4e, 16'h9c4e, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4e, 16'h9c2d, 16'h9c4e, 16'h9c4f, 16'h9c4f, 16'h9c2e, 16'h7b2a, 16'h41a5, 16'h3144, 16'h2944, 16'h213, 16'h820, 16'h861, 16'h861, 16'h020, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2923, 16'h2923, 16'h6a86, 16'h6a86, 16'h5a47, 16'h5a47, 16'h5a47, 16'h5a47, 16'h5a47, 16'h5a47, 16'h5a47, 16'h5a47, 16'h6267, 16'h6aa9, 16'h94d, 16'h7b4a, 16'h41c5, 16'h1081, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h840, 16'h3144, 16'h9c4f, 16'hacd1, 16'hacd0, 16'hacb0, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha46f, 16'ha470, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4e, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9ce, 16'h9ce, 16'h9cd, 16'h94d, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h8bcd, 16'h93cd, 16'h93cd, 16'h8bcd, 16'h8bcd, 16'h8bcd, 16'h8bcc, 16'h8bcc, 16'h8bac, 16'h8bac, 16'h8bac, 16'h8bac, 16'h8bac, 16'h8bac, 16'h8bac, 16'h8b8d, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h838b, 16'h838b, 16'h838b, 16'h836b, 16'h836b, 16'h7b4a, 16'h49e6, 16'h212, 16'h20e1, 16'h20c2, 16'h20c1, 16'h18c1, 16'h820, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h7b4b, 16'h834b, 16'h836b, 16'h836b, 16'h836c, 16'h836c, 16'h836b, 16'h7b4b, 16'h836c, 16'h836c, 16'h836c, 16'h838c, 16'h73a, 16'h62a9, 16'h62a9, 16'h73a, 16'h836c, 16'h8bad, 16'h8bad, 16'h8bad, 16'h8bad, 16'h93ee, 16'h8bcd, 16'h942e, 16'h9c2e, 16'h9c4e, 16'h9c4e, 16'h9c4f, 16'h9c4e, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4e, 16'h9c4e, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4e, 16'h7b2a, 16'h41a5, 16'h3144, 16'h2944, 16'h213, 16'h820, 16'h861, 16'h861, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h020, 16'h00, 16'h00, 16'h18c2, 16'h293, 16'h72a6, 16'h6a86, 16'h5a46, 16'h5a47, 16'h5a47, 16'h5a47, 16'h5a47, 16'h5a47, 16'h5a47, 16'h5a47, 16'h6267, 16'h6aa9, 16'h93ed, 16'h7b4a, 16'h41c5, 16'h1081, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h840, 16'h3124, 16'ha44f, 16'hacd1, 16'hacd0, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha46f, 16'ha470, 16'ha450, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9ce, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9ce, 16'h9c2e, 16'h9ce, 16'h9ce, 16'h94d, 16'h94e, 16'h93ee, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93cd, 16'h93ed, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h8bcd, 16'h8bcd, 16'h8bcd, 16'h8bcc, 16'h8bcc, 16'h8bad, 16'h8bad, 16'h8bad, 16'h8bac, 16'h8bad, 16'h8bac, 16'h8bac, 16'h8bac, 16'h8bac, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8b, 16'h838c, 16'h836c, 16'h838c, 16'h836c, 16'h836b, 16'h7b4b, 16'h49e6, 16'h20e2, 16'h20e2, 16'h20e2, 16'h20e1, 16'h18a1, 16'h820, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h7b4b, 16'h834c, 16'h836b, 16'h7b4b, 16'h7b2b, 16'h7b4b, 16'h7b4b, 16'h7b4b, 16'h836c, 16'h836c, 16'h7b6b, 16'h7b8c, 16'h732a, 16'h62a9, 16'h62a9, 16'h72ea, 16'h7b4c, 16'h83ad, 16'h8bcd, 16'h8bad, 16'h8bad, 16'h8bed, 16'h8bed, 16'h942e, 16'h942e, 16'h9c4e, 16'h9c4e, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c6e, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c50, 16'h9c4f, 16'h7b2a, 16'h49c5, 16'h3164, 16'h3144, 16'h213, 16'h840, 16'h861, 16'h1061, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h00, 16'h00, 16'h860, 16'h20e2, 16'h72a6, 16'h6a87, 16'h5a47, 16'h5a47, 16'h5a47, 16'h5a47, 16'h5a47, 16'h5a47, 16'h5a47, 16'h5a47, 16'h6267, 16'h6aa9, 16'h93cd, 16'h7b2a, 16'h41c5, 16'h1081, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h820, 16'h840, 16'h3144, 16'ha44f, 16'hacb1, 16'hacd0, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha470, 16'ha450, 16'ha450, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c2f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9ce, 16'h9ce, 16'h9ce, 16'h9c2e, 16'h9ce, 16'h9ce, 16'h9ce, 16'h94e, 16'h94d, 16'h94e, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93cd, 16'h93cd, 16'h93cd, 16'h8bcd, 16'h93cd, 16'h8bcd, 16'h8bcd, 16'h8bcd, 16'h8bcd, 16'h8bcc, 16'h8bac, 16'h8bac, 16'h8bac, 16'h8bac, 16'h8bac, 16'h8bad, 16'h8bad, 16'h8b8d, 16'h8bac, 16'h8bac, 16'h8bac, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h838c, 16'h838c, 16'h836c, 16'h838c, 16'h836c, 16'h836c, 16'h7b4a, 16'h49e6, 16'h20e2, 16'h20e1, 16'h20e2, 16'h20e1, 16'h18a1, 16'h820, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h7b6b, 16'h834b, 16'h7b4b, 16'h732b, 16'h73a, 16'h72ea, 16'h7b2b, 16'h7b4b, 16'h7b6b, 16'h7b6b, 16'h7b6b, 16'h7b6c, 16'h732a, 16'h62a9, 16'h62a9, 16'h72ea, 16'h7b6c, 16'h83ac, 16'h8bad, 16'h8bac, 16'h8bad, 16'h8bed, 16'h93ed, 16'h942e, 16'h942e, 16'h9c2e, 16'h9c4e, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c6f, 16'h9c6f, 16'h9c6f, 16'h9c6f, 16'h9c70, 16'h9c4f, 16'h7b4b, 16'h49c6, 16'h3164, 16'h3164, 16'h2924, 16'h841, 16'h841, 16'h1081, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h00, 16'h1081, 16'h18a1, 16'h6a85, 16'h6a87, 16'h5a47, 16'h5a47, 16'h5a47, 16'h5a46, 16'h5a47, 16'h5a47, 16'h5a47, 16'h5a47, 16'h6267, 16'h6aa9, 16'h93cc, 16'h7ba, 16'h49c5, 16'h1081, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h840, 16'h840, 16'h3144, 16'ha44f, 16'hacb1, 16'hacb1, 16'hacd0, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha450, 16'ha450, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9ce, 16'h9ce, 16'h9ce, 16'h9ce, 16'h94e, 16'h9ce, 16'h94e, 16'h94d, 16'h94d, 16'h94e, 16'h93ee, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93cd, 16'h8bed, 16'h93cd, 16'h8bcd, 16'h8bcd, 16'h8bcd, 16'h8bcd, 16'h8bcd, 16'h8bcd, 16'h8bad, 16'h8bad, 16'h8bad, 16'h8bad, 16'h8bac, 16'h8bac, 16'h8bac, 16'h8bac, 16'h8bac, 16'h8bac, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8b, 16'h8b8b, 16'h8b8b, 16'h838b, 16'h836b, 16'h836c, 16'h836b, 16'h7b4a, 16'h49e6, 16'h20e2, 16'h20e1, 16'h20e1, 16'h20e1, 16'h18c1, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h7b4b, 16'h7b4b, 16'h7b2b, 16'h72ea, 16'h72ea, 16'h72ea, 16'h7b2b, 16'h7b2b, 16'h7b4b, 16'h7b6b, 16'h7b6b, 16'h7b6c, 16'h7b2b, 16'h6ac9, 16'h6aea, 16'h7b4b, 16'h838c, 16'h83ac, 16'h8bac, 16'h8bac, 16'h8bcd, 16'h93ed, 16'h94d, 16'h94d, 16'h942e, 16'h9c2e, 16'h9c4e, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c6f, 16'h9c6f, 16'h9c6f, 16'h9c6f, 16'ha46f, 16'ha470, 16'ha470, 16'ha46f, 16'h836b, 16'h49c6, 16'h3164, 16'h3164, 16'h2924, 16'h841, 16'h841, 16'h1081, 16'h020, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h00, 16'h1081, 16'h20c2, 16'h6a66, 16'h6a87, 16'h5a47, 16'h5a47, 16'h5a47, 16'h5a46, 16'h5a46, 16'h5a47, 16'h5a47, 16'h5a47, 16'h5a47, 16'h6aa9, 16'h93cc, 16'h7ba, 16'h49c5, 16'h1081, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h00, 16'h020, 16'h020, 16'h020, 16'h040, 16'h840, 16'h3143, 16'ha44f, 16'hacb1, 16'hacb1, 16'hacb0, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha470, 16'ha46f, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9ce, 16'h9ce, 16'h9ce, 16'h9cd, 16'h9ce, 16'h9ce, 16'h94e, 16'h94d, 16'h94d, 16'h94d, 16'h94d, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93cd, 16'h93cd, 16'h8bcd, 16'h8bcd, 16'h8bcd, 16'h8bcd, 16'h8bcd, 16'h8bcd, 16'h8bcd, 16'h8bad, 16'h8bad, 16'h8bad, 16'h8bad, 16'h8bad, 16'h8bac, 16'h8bac, 16'h8bac, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8b, 16'h8b8c, 16'h836c, 16'h836b, 16'h836b, 16'h836b, 16'h7b4a, 16'h49e5, 16'h20e1, 16'h20e1, 16'h20c1, 16'h20c1, 16'h18c1, 16'h820, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h7b4b, 16'h7b4b, 16'h7b2a, 16'h73a, 16'h7b2b, 16'h7b2b, 16'h732a, 16'h7b2a, 16'h7b4b, 16'h7b6b, 16'h7b6b, 16'h7b6b, 16'h7b6b, 16'h7b6b, 16'h836c, 16'h838b, 16'h83ac, 16'h83ac, 16'h8bcc, 16'h8bcd, 16'h8bed, 16'h8cd, 16'h94d, 16'h94e, 16'h942e, 16'h9c2e, 16'h9c4e, 16'h9c4f, 16'h9c4f, 16'h9c6f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha470, 16'ha490, 16'ha490, 16'ha490, 16'h838b, 16'h49c5, 16'h3164, 16'h3184, 16'h2944, 16'h841, 16'h841, 16'h10a1, 16'h020, 16'h00, 16'h00, 16'h020, 16'h820, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h841, 16'h2923, 16'h292, 16'h6a66, 16'h6a87, 16'h5a47, 16'h5a47, 16'h5a47, 16'h5a47, 16'h5a47, 16'h5a47, 16'h5a47, 16'h5a47, 16'h5a47, 16'h6aa8, 16'h93cc, 16'h732a, 16'h41c5, 16'h1081, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h020, 16'h00, 16'h020, 16'h020, 16'h020, 16'h040, 16'h840, 16'h3143, 16'ha44f, 16'hacb1, 16'hacb1, 16'hacd0, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h94e, 16'h9ce, 16'h9ce, 16'h94e, 16'h94e, 16'h94d, 16'h94d, 16'h94d, 16'h94d, 16'h94d, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h8bcd, 16'h8bcd, 16'h8bcd, 16'h8bcd, 16'h8bcd, 16'h8bad, 16'h8bad, 16'h8bad, 16'h8bac, 16'h8bad, 16'h8bac, 16'h8bac, 16'h8bac, 16'h8b8c, 16'h8b8c, 16'h8b8d, 16'h8b8d, 16'h8b8c, 16'h8b8c, 16'h838c, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h838b, 16'h838b, 16'h836c, 16'h836c, 16'h836c, 16'h836b, 16'h7b4b, 16'h49e6, 16'h20e1, 16'h20c1, 16'h20c1, 16'h20c1, 16'h18c1, 16'h820, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h7b2a, 16'h7b2a, 16'h73a, 16'h73a, 16'h73a, 16'h73a, 16'h73a, 16'h7b2a, 16'h7b4a, 16'h7b4b, 16'h7b4b, 16'h7b4b, 16'h7b6b, 16'h836b, 16'h838b, 16'h838b, 16'h83ac, 16'h8bac, 16'h8bcc, 16'h8bed, 16'h8bed, 16'h93ed, 16'h94d, 16'h94d, 16'h942e, 16'h9c2e, 16'h9c4e, 16'h9c4e, 16'h9c4f, 16'h9c6f, 16'h9c6f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h94e, 16'h8bcd, 16'h6ac9, 16'h41c6, 16'h3185, 16'h3985, 16'h3164, 16'h861, 16'h841, 16'h10a1, 16'h020, 16'h00, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h00, 16'h020, 16'h00, 16'h00, 16'h00, 16'h820, 16'h1081, 16'h18c1, 16'h861, 16'h020, 16'h020, 16'h020, 16'h020, 16'h1061, 16'h5a47, 16'h6267, 16'h838, 16'h6a87, 16'h5a47, 16'h5a47, 16'h5a47, 16'h5a46, 16'h5a46, 16'h5a27, 16'h5a47, 16'h5a47, 16'h6247, 16'h6aa8, 16'h93cc, 16'h732a, 16'h41c5, 16'h1081, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h040, 16'h3144, 16'ha44f, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha470, 16'ha46f, 16'ha470, 16'ha470, 16'ha46f, 16'ha46f, 16'ha450, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h9c4e, 16'h9c2e, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9ce, 16'h9c2e, 16'h9ce, 16'h94e, 16'h94e, 16'h9cd, 16'h94d, 16'h94d, 16'h94d, 16'h94d, 16'h94d, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h8bcc, 16'h8bac, 16'h8bac, 16'h8bac, 16'h8bac, 16'h8bad, 16'h8bac, 16'h8bac, 16'h8bac, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h838c, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h838c, 16'h838b, 16'h836c, 16'h836b, 16'h836b, 16'h836b, 16'h7b4a, 16'h49e5, 16'h20e1, 16'h20c1, 16'h20c1, 16'h20c1, 16'h18a1, 16'h820, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h73a, 16'h73a, 16'h73a, 16'h73a, 16'h732a, 16'h732a, 16'h7b2b, 16'h7b4b, 16'h7b4b, 16'h7b4b, 16'h7b4b, 16'h7b4b, 16'h7b6b, 16'h7b6a, 16'h838b, 16'h838b, 16'h83ab, 16'h83ac, 16'h8bcc, 16'h8bcd, 16'h8bed, 16'h94d, 16'h94d, 16'h94d, 16'h942d, 16'h942e, 16'h9c4d, 16'h9c4e, 16'h942e, 16'h94d, 16'h83cd, 16'h7b6c, 16'h6aea, 16'h5a88, 16'h4a7, 16'h3185, 16'h213, 16'h18a2, 16'h20c3, 16'h41a5, 16'h39a5, 16'h39a5, 16'h3184, 16'h861, 16'h841, 16'h10a2, 16'h020, 16'h00, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h1061, 16'h2923, 16'h2923, 16'h1081, 16'h020, 16'h020, 16'h040, 16'h020, 16'h1081, 16'h5a67, 16'h836a, 16'ha4b, 16'h6a87, 16'h5a47, 16'h5a27, 16'h5a27, 16'h5a46, 16'h5a46, 16'h5a47, 16'h5a47, 16'h5a47, 16'h5a47, 16'h6aa8, 16'h8bcc, 16'h732a, 16'h41c5, 16'h1081, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h00, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h040, 16'h3144, 16'h9c4f, 16'hacd0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'ha490, 16'ha48f, 16'ha470, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c2f, 16'h9c4f, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9ce, 16'h9c2e, 16'h9c2e, 16'h9ce, 16'h9ce, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94d, 16'h94d, 16'h94d, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h8bad, 16'h8bad, 16'h8bac, 16'h8bac, 16'h8bad, 16'h8bad, 16'h8bac, 16'h8bac, 16'h8bac, 16'h8bac, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h838c, 16'h8b8c, 16'h8b8c, 16'h838c, 16'h838b, 16'h8b8b, 16'h838c, 16'h838b, 16'h836b, 16'h836b, 16'h7b2a, 16'h49e5, 16'h20e1, 16'h20c1, 16'h20c1, 16'h20c1, 16'h18a1, 16'h820, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h73a, 16'h73a, 16'h73a, 16'h73a, 16'h732a, 16'h732a, 16'h732a, 16'h7b2a, 16'h7b4a, 16'h7b4a, 16'h7b4a, 16'h7b4a, 16'h7b4a, 16'h7b6a, 16'h836b, 16'h838b, 16'h838b, 16'h83ac, 16'h8bac, 16'h8bcc, 16'h8bcd, 16'h8bed, 16'h94d, 16'h94d, 16'h94e, 16'h942e, 16'h942e, 16'h8bcd, 16'h4a7, 16'h2944, 16'h18e3, 16'h1082, 16'h861, 16'h840, 16'h040, 16'h020, 16'h020, 16'h020, 16'h1081, 16'h41a5, 16'h41a5, 16'h41a6, 16'h3185, 16'h861, 16'h841, 16'h18c2, 16'h020, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h00, 16'h00, 16'h00, 16'h1061, 16'h2943, 16'h2923, 16'h1081, 16'h020, 16'h020, 16'h040, 16'h020, 16'h18a1, 16'h6ac8, 16'h834a, 16'ha42b, 16'h6a87, 16'h5a47, 16'h5a46, 16'h5a46, 16'h5a46, 16'h5a46, 16'h5a47, 16'h5a47, 16'h5a47, 16'h6267, 16'h6aa8, 16'h8bcc, 16'h732a, 16'h41c5, 16'h1081, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h020, 16'h040, 16'h3144, 16'h9c6f, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9ce, 16'h9c2e, 16'h9ce, 16'h9ce, 16'h9ce, 16'h9ce, 16'h94e, 16'h94e, 16'h94e, 16'h94d, 16'h94d, 16'h94d, 16'h94d, 16'h94d, 16'h94d, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h8bcd, 16'h8bcd, 16'h8bcd, 16'h8bcd, 16'h8bcc, 16'h8bad, 16'h8bad, 16'h8bac, 16'h8bac, 16'h8bac, 16'h8bac, 16'h8bac, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h838c, 16'h838c, 16'h838c, 16'h8b8c, 16'h8b8c, 16'h838b, 16'h838b, 16'h836c, 16'h836b, 16'h836c, 16'h836b, 16'h7b2b, 16'h49c5, 16'h20e1, 16'h20c1, 16'h20c1, 16'h20e0, 16'h18c1, 16'h820, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h739, 16'h73a, 16'h73a, 16'h73a, 16'h73a, 16'h73a, 16'h732a, 16'h732a, 16'h7b2a, 16'h7b2a, 16'h7b2b, 16'h7b4a, 16'h7b4a, 16'h7b6b, 16'h7b6b, 16'h836b, 16'h838b, 16'h83ac, 16'h83ac, 16'h8bcc, 16'h8bcd, 16'h8bec, 16'h93ed, 16'h94d, 16'h94e, 16'h942e, 16'h942e, 16'h838c, 16'h20e2, 16'h840, 16'h040, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h1081, 16'h39a5, 16'h41c5, 16'h41c5, 16'h31a5, 16'h1081, 16'h841, 16'h18c2, 16'h020, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h00, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h00, 16'h00, 16'h00, 16'h1061, 16'h2943, 16'h3143, 16'h10a1, 16'h020, 16'h020, 16'h020, 16'h840, 16'h18a1, 16'h6287, 16'h834a, 16'h9beb, 16'h6a66, 16'h5a26, 16'h5a27, 16'h5a47, 16'h5a46, 16'h5a46, 16'h5a27, 16'h5a47, 16'h5a46, 16'h6267, 16'h6aa8, 16'h8bcc, 16'h7b2a, 16'h49c5, 16'h1081, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h3144, 16'ha46f, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9ce, 16'h9ce, 16'h9ce, 16'h9ce, 16'h9ce, 16'h9ce, 16'h9ce, 16'h94e, 16'h94e, 16'h94d, 16'h94e, 16'h93ee, 16'h94d, 16'h94d, 16'h93ed, 16'h94d, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h8bcd, 16'h8bcd, 16'h8bcd, 16'h8bcd, 16'h8bad, 16'h8bac, 16'h8bac, 16'h8bad, 16'h8bad, 16'h8bac, 16'h8bac, 16'h8bac, 16'h8b8c, 16'h8b8d, 16'h8b8d, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h838c, 16'h838c, 16'h838c, 16'h838c, 16'h8b8c, 16'h8b8c, 16'h838b, 16'h838b, 16'h836b, 16'h836b, 16'h836b, 16'h836b, 16'h7b2b, 16'h49c5, 16'h20e2, 16'h20c1, 16'h18c1, 16'h18c1, 16'h18a1, 16'h820, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h6ae9, 16'h6ba, 16'h6ba, 16'h6ba, 16'h73a, 16'h73a, 16'h73a, 16'h73a, 16'h7b2a, 16'h7b2a, 16'h7b2b, 16'h7b4a, 16'h7b4a, 16'h7b4b, 16'h7b6b, 16'h836b, 16'h838b, 16'h83ab, 16'h83ac, 16'h8bac, 16'h8bcc, 16'h8bcd, 16'h93ed, 16'h94d, 16'h94d, 16'h94d, 16'h942e, 16'h838b, 16'h192, 16'h040, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h1081, 16'h39a5, 16'h41c6, 16'h41c6, 16'h39c6, 16'h10a2, 16'h841, 16'h18c2, 16'h020, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h00, 16'h020, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h00, 16'h00, 16'h00, 16'h1061, 16'h2123, 16'h213, 16'h1081, 16'h020, 16'h020, 16'h020, 16'h020, 16'h213, 16'h5a66, 16'h5a47, 16'h8328, 16'h6a86, 16'h5225, 16'h5a26, 16'h5a47, 16'h5a47, 16'h5a46, 16'h5a46, 16'h5a46, 16'h5a46, 16'h6267, 16'h6aa8, 16'h8bcc, 16'h7b2a, 16'h49c5, 16'h1081, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h3144, 16'h9c4f, 16'hacb0, 16'hacd0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'hacb1, 16'hb4d1, 16'hacb0, 16'ha490, 16'ha46f, 16'ha470, 16'ha470, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9ce, 16'h9ce, 16'h9c2e, 16'h9ce, 16'h9ce, 16'h9ce, 16'h9ce, 16'h94e, 16'h94e, 16'h94e, 16'h94d, 16'h94d, 16'h93ed, 16'h94d, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h8bcd, 16'h8bcd, 16'h8bcd, 16'h8bcd, 16'h8bcd, 16'h8bad, 16'h8bad, 16'h8bac, 16'h8bad, 16'h8bac, 16'h8bad, 16'h8bac, 16'h8bac, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h836c, 16'h838c, 16'h838c, 16'h8b6c, 16'h836c, 16'h838b, 16'h838b, 16'h836b, 16'h836b, 16'h838b, 16'h836b, 16'h7b2a, 16'h41e5, 16'h20e1, 16'h20c1, 16'h18c1, 16'h18c1, 16'h18a0, 16'h820, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h6ae9, 16'h6ae9, 16'h6aea, 16'h739, 16'h739, 16'h73a, 16'h73a, 16'h73a, 16'h73a, 16'h732a, 16'h7b2a, 16'h7b4a, 16'h7b4a, 16'h7b4a, 16'h7b6a, 16'h836b, 16'h838b, 16'h838b, 16'h83ac, 16'h8bac, 16'h8bcc, 16'h8bcc, 16'h8bed, 16'h93ed, 16'h94d, 16'h94d, 16'h942d, 16'h7b8b, 16'h212, 16'h040, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h1081, 16'h39a5, 16'h49e6, 16'h41e6, 16'h41c6, 16'h10a2, 16'h841, 16'h18c2, 16'h020, 16'h00, 16'h00, 16'h020, 16'h020, 16'h00, 16'h00, 16'h020, 16'h020, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h841, 16'h820, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h3164, 16'h8bca, 16'h93eb, 16'h93a9, 16'h6aa7, 16'h5a46, 16'h5a46, 16'h5a47, 16'h5a46, 16'h5a46, 16'h5a46, 16'h5a46, 16'h5a46, 16'h6267, 16'h6aa8, 16'h8bac, 16'h7b2a, 16'h41c5, 16'h1081, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h3144, 16'h9c6f, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'hacb1, 16'hb4d1, 16'hb4d1, 16'hac90, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha46f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9ce, 16'h9ce, 16'h9ce, 16'h9ce, 16'h94d, 16'h94d, 16'h94d, 16'h94e, 16'h94e, 16'h94d, 16'h94d, 16'h93ed, 16'h93ed, 16'h94d, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93cd, 16'h93cd, 16'h8bcd, 16'h8bcd, 16'h93cd, 16'h8bcd, 16'h8bcd, 16'h8bcd, 16'h8bcd, 16'h8bcd, 16'h8bad, 16'h8bad, 16'h8bac, 16'h8bac, 16'h8bad, 16'h8bad, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h838c, 16'h838b, 16'h8b8c, 16'h836c, 16'h838b, 16'h838b, 16'h836b, 16'h836b, 16'h836b, 16'h836b, 16'h7b2a, 16'h49e5, 16'h20e1, 16'h20c1, 16'h18c1, 16'h18e1, 16'h18c0, 16'h820, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h6ae9, 16'h6ae9, 16'h6ae9, 16'h72ea, 16'h739, 16'h6ba, 16'h73a, 16'h73a, 16'h73a, 16'h732a, 16'h732a, 16'h732a, 16'h7b2a, 16'h7b4a, 16'h7b4a, 16'h836a, 16'h838b, 16'h838b, 16'h838b, 16'h8bac, 16'h8bcc, 16'h8bcc, 16'h8bcd, 16'h8bed, 16'h93ed, 16'h94d, 16'h94d, 16'h7b8b, 16'h212, 16'h840, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h040, 16'h040, 16'h020, 16'h861, 16'h39a5, 16'h4a7, 16'h41e6, 16'h41c6, 16'h18a2, 16'h841, 16'h18c2, 16'h020, 16'h00, 16'h00, 16'h00, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h840, 16'h3964, 16'h8349, 16'ha44d, 16'ha42c, 16'h6aa7, 16'h5a46, 16'h5a46, 16'h5a47, 16'h5a46, 16'h5a46, 16'h5a46, 16'h5a46, 16'h5a46, 16'h6247, 16'h6aa8, 16'h8bcc, 16'h7b29, 16'h41c4, 16'h1081, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h3144, 16'h9c6f, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'hac90, 16'hacb0, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9ce, 16'h9ce, 16'h9ce, 16'h94e, 16'h94e, 16'h94d, 16'h94d, 16'h94e, 16'h94e, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93cd, 16'h93cd, 16'h93cd, 16'h8bcd, 16'h8bcd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h8bcd, 16'h8bcd, 16'h8bad, 16'h8bad, 16'h8bac, 16'h8bac, 16'h8bad, 16'h8bad, 16'h8bac, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b6c, 16'h838c, 16'h8b8b, 16'h8b8b, 16'h836b, 16'h838b, 16'h836c, 16'h836c, 16'h836b, 16'h836b, 16'h7b2a, 16'h49e5, 16'h20e1, 16'h20c1, 16'h20c1, 16'h18c1, 16'h18a1, 16'h820, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h6ae9, 16'h6ae9, 16'h6ae9, 16'h6aea, 16'h6aea, 16'h6ba, 16'h6ba, 16'h73a, 16'h73a, 16'h732a, 16'h732a, 16'h732a, 16'h7b2a, 16'h7b2a, 16'h7b4a, 16'h7b4b, 16'h836b, 16'h838b, 16'h838b, 16'h83ab, 16'h8bac, 16'h8bac, 16'h8bcd, 16'h8bec, 16'h93ed, 16'h94d, 16'h94d, 16'h7b8b, 16'h212, 16'h040, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h040, 16'h040, 16'h020, 16'h861, 16'h39a5, 16'h4a27, 16'h4a7, 16'h41e6, 16'h18c2, 16'h841, 16'h18e3, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h840, 16'h525, 16'h8baa, 16'h9cc, 16'ha4b, 16'h6aa7, 16'h5a46, 16'h5a46, 16'h5a46, 16'h5a27, 16'h5a47, 16'h5a46, 16'h5a46, 16'h5a46, 16'h6267, 16'h6aa8, 16'h8bac, 16'h7b4a, 16'h41c4, 16'h1081, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h3144, 16'ha46f, 16'hacd0, 16'hacd0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha46f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c2e, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9ce, 16'h9ce, 16'h9ce, 16'h94e, 16'h94e, 16'h94d, 16'h94e, 16'h94d, 16'h94e, 16'h94d, 16'h94d, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93cd, 16'h93cd, 16'h93cd, 16'h8bcd, 16'h8bcd, 16'h93cd, 16'h8bcd, 16'h8bad, 16'h8bcd, 16'h8bcd, 16'h8bad, 16'h8bad, 16'h8bac, 16'h8bac, 16'h8bac, 16'h8b8c, 16'h8bac, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8b, 16'h8b6c, 16'h836c, 16'h838c, 16'h838b, 16'h836c, 16'h836b, 16'h836b, 16'h836b, 16'h7b2b, 16'h41c5, 16'h20e1, 16'h18c1, 16'h20c1, 16'h20c1, 16'h10a0, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h6ae9, 16'h6ae9, 16'h6ae9, 16'h6ac9, 16'h6ae9, 16'h6aea, 16'h6aea, 16'h72e9, 16'h73a, 16'h73a, 16'h73a, 16'h732a, 16'h732a, 16'h7b2a, 16'h7b4a, 16'h7b4a, 16'h7b6a, 16'h7b6a, 16'h838b, 16'h838b, 16'h83ab, 16'h8bac, 16'h8bcc, 16'h8bcc, 16'h8bcd, 16'h8bed, 16'h8cc, 16'h7b8a, 16'h2122, 16'h040, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h861, 16'h39a5, 16'h5227, 16'h4a7, 16'h4a7, 16'h18e2, 16'h841, 16'h18e2, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h840, 16'h18a1, 16'h5225, 16'h8349, 16'h93cc, 16'ha4c, 16'h6aa7, 16'h5a46, 16'h5a46, 16'h5a26, 16'h5227, 16'h5a46, 16'h5a46, 16'h5a46, 16'h5a46, 16'h5a66, 16'h6aa8, 16'h8bcc, 16'h7b49, 16'h41c4, 16'h1081, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h3164, 16'ha46f, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c2e, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9ce, 16'h9ce, 16'h9c2e, 16'h9ce, 16'h9ce, 16'h94e, 16'h94e, 16'h94e, 16'h94d, 16'h94d, 16'h94d, 16'h93ee, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h8bcd, 16'h8bcd, 16'h8bcd, 16'h8bcd, 16'h8bcd, 16'h8bad, 16'h8bac, 16'h8bac, 16'h8bac, 16'h8bac, 16'h8bac, 16'h8bac, 16'h8b8c, 16'h8bac, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b6c, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8b, 16'h8b6c, 16'h836c, 16'h836b, 16'h836b, 16'h836b, 16'h836b, 16'h836b, 16'h836b, 16'h7b2a, 16'h41c5, 16'h20e2, 16'h18c1, 16'h20c1, 16'h20c1, 16'h18a0, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h6ac9, 16'h6ac9, 16'h6ae9, 16'h6ae9, 16'h6ae9, 16'h6ae9, 16'h6ae9, 16'h6ae9, 16'h6aea, 16'h6b9, 16'h6b9, 16'h73a, 16'h732a, 16'h732a, 16'h7b2a, 16'h7b4a, 16'h7b4a, 16'h7b6a, 16'h7b6b, 16'h836b, 16'h838b, 16'h83ab, 16'h8bac, 16'h8bcc, 16'h8bcc, 16'h8bcc, 16'h8bec, 16'h7b6a, 16'h2122, 16'h040, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h861, 16'h3985, 16'h5247, 16'h4a27, 16'h4a7, 16'h20e3, 16'h841, 16'h20e2, 16'h820, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h860, 16'h1081, 16'h20c1, 16'h5a46, 16'h7b28, 16'h8baa, 16'h9bea, 16'h72a7, 16'h5a26, 16'h5a27, 16'h5a26, 16'h5a26, 16'h5a26, 16'h5a46, 16'h5a46, 16'h5a46, 16'h5a67, 16'h6aa8, 16'h8bac, 16'h7b2a, 16'h41c5, 16'h1081, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h3164, 16'ha46f, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha470, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9ce, 16'h9ce, 16'h9ce, 16'h9ce, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94d, 16'h94d, 16'h94d, 16'h94d, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93cd, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93cd, 16'h93cd, 16'h93cd, 16'h8bad, 16'h8bad, 16'h8bad, 16'h8bad, 16'h8bcd, 16'h8bad, 16'h8bad, 16'h8bac, 16'h8bad, 16'h8bad, 16'h8bac, 16'h8bac, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8b, 16'h8b8b, 16'h8b8b, 16'h8b8b, 16'h836c, 16'h838b, 16'h836b, 16'h836b, 16'h836c, 16'h836b, 16'h836b, 16'h836b, 16'h7b2a, 16'h49c5, 16'h20e1, 16'h18c1, 16'h18c1, 16'h18c0, 16'h10a0, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h6ac8, 16'h6ac9, 16'h6ac9, 16'h6ac9, 16'h6ae9, 16'h6ac9, 16'h6ae9, 16'h6ae9, 16'h6ae9, 16'h6b9, 16'h6b9, 16'h6b9, 16'h739, 16'h73a, 16'h732a, 16'h7b2a, 16'h7b4a, 16'h7b4b, 16'h7b6b, 16'h836b, 16'h838b, 16'h838b, 16'h838b, 16'h83ab, 16'h8bac, 16'h8bac, 16'h8bcc, 16'h7329, 16'h212, 16'h840, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h861, 16'h3985, 16'h5248, 16'h5227, 16'h4a26, 16'h213, 16'h820, 16'h212, 16'h820, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h00, 16'h00, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h840, 16'h860, 16'h1080, 16'h1080, 16'h20c1, 16'h72e8, 16'h93ca, 16'hac8e, 16'ha42c, 16'h6aa6, 16'h5a46, 16'h5a26, 16'h5a26, 16'h5a26, 16'h5a26, 16'h5a26, 16'h5a27, 16'h5a47, 16'h5a67, 16'h6aa8, 16'h8bab, 16'h7b4a, 16'h41c5, 16'h1081, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h820, 16'h3164, 16'ha46f, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9ce, 16'h9ce, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h93ee, 16'h94d, 16'h93ed, 16'h93ed, 16'h93ee, 16'h93ed, 16'h93ed, 16'h93ee, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h8bad, 16'h8bad, 16'h8bad, 16'h8bad, 16'h8bad, 16'h8bad, 16'h8bad, 16'h8bad, 16'h8bad, 16'h8bad, 16'h8bac, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8b, 16'h838b, 16'h838b, 16'h8b6c, 16'h836b, 16'h836b, 16'h836b, 16'h836c, 16'h836b, 16'h836b, 16'h834c, 16'h7b2b, 16'h49c5, 16'h20e1, 16'h18c1, 16'h18c1, 16'h18c1, 16'h10a1, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h62a8, 16'h62c8, 16'h62c9, 16'h62c8, 16'h6ae8, 16'h6ac9, 16'h6ae9, 16'h6ae9, 16'h6ae9, 16'h6ae9, 16'h6aea, 16'h6aea, 16'h6ba, 16'h73a, 16'h73a, 16'h7329, 16'h7b4a, 16'h7b4a, 16'h7b4b, 16'h836b, 16'h836b, 16'h838b, 16'h838b, 16'h838b, 16'h83ab, 16'h8bac, 16'h838b, 16'h5a67, 16'h18e2, 16'h040, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h861, 16'h39a5, 16'h5a68, 16'h5227, 16'h4a27, 16'h213, 16'h820, 16'h213, 16'h840, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h00, 16'h00, 16'h00, 16'h020, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h020, 16'h040, 16'h860, 16'h860, 16'h1080, 16'h1080, 16'h18c1, 16'h62a7, 16'h8b8a, 16'h8baa, 16'h9389, 16'h6aa7, 16'h5a47, 16'h5a46, 16'h5a26, 16'h5a46, 16'h5a27, 16'h5a27, 16'h5a27, 16'h5a47, 16'h5a66, 16'h6aa8, 16'h8bab, 16'h7b49, 16'h41e4, 16'h1081, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h840, 16'h3164, 16'ha46f, 16'hacd1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac8f, 16'ha490, 16'ha490, 16'ha490, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha470, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9ce, 16'h94e, 16'h9ce, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h93ee, 16'h94e, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93cd, 16'h93cd, 16'h8bcd, 16'h93cd, 16'h8bcd, 16'h93cc, 16'h8bac, 16'h8bac, 16'h8bad, 16'h8bad, 16'h8bad, 16'h8bad, 16'h8bac, 16'h8bac, 16'h8bac, 16'h8bac, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h838c, 16'h838b, 16'h838b, 16'h836b, 16'h836c, 16'h836b, 16'h836c, 16'h836b, 16'h836b, 16'h836b, 16'h7b2a, 16'h41c5, 16'h20e1, 16'h18c1, 16'h18c1, 16'h18e0, 16'h10a0, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h62a8, 16'h62a8, 16'h62a8, 16'h62c8, 16'h6ac8, 16'h6ac9, 16'h6ac9, 16'h6ae9, 16'h6ae9, 16'h6ae9, 16'h6aea, 16'h6aea, 16'h6b9, 16'h72ea, 16'h73a, 16'h7329, 16'h732a, 16'h732a, 16'h7b4a, 16'h7b4a, 16'h7b6a, 16'h836b, 16'h836b, 16'h838b, 16'h838b, 16'h838b, 16'h6ae9, 16'h41e4, 16'h10c1, 16'h040, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h841, 16'h39a5, 16'h5a89, 16'h5a47, 16'h5247, 16'h2123, 16'h820, 16'h213, 16'h840, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h040, 16'h860, 16'h880, 16'h880, 16'h880, 16'h18a1, 16'h6267, 16'h72c8, 16'h7b9, 16'h93ca, 16'h72a7, 16'h5a26, 16'h5a46, 16'h5a26, 16'h5a26, 16'h5a27, 16'h5a26, 16'h5a46, 16'h5a46, 16'h5a67, 16'h6aa8, 16'h8bac, 16'h7b4a, 16'h41e5, 16'h1081, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h040, 16'h3164, 16'ha46f, 16'hacd0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha48f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c4f, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9ce, 16'h9ce, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94d, 16'h94d, 16'h94d, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h8bcd, 16'h8bcd, 16'h8bad, 16'h8bac, 16'h8bad, 16'h8bad, 16'h8bac, 16'h8bad, 16'h8bad, 16'h8bac, 16'h8bac, 16'h8bac, 16'h8bac, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h838c, 16'h838c, 16'h8b8c, 16'h8b8c, 16'h8b8b, 16'h8b8c, 16'h838c, 16'h838c, 16'h838c, 16'h838c, 16'h836c, 16'h836b, 16'h836b, 16'h836c, 16'h836b, 16'h836b, 16'h836b, 16'h7b2a, 16'h41c5, 16'h20e1, 16'h20e1, 16'h18c1, 16'h18e1, 16'h10a0, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h62a8, 16'h62a8, 16'h62a8, 16'h62a8, 16'h62a8, 16'h6aa9, 16'h6ac9, 16'h6ac9, 16'h6ac9, 16'h6ac9, 16'h6ac9, 16'h6ae9, 16'h6ae9, 16'h72e9, 16'h6aea, 16'h739, 16'h73a, 16'h732a, 16'h7b2a, 16'h7b4a, 16'h7b4a, 16'h7b4b, 16'h7b4b, 16'h836b, 16'h7b6b, 16'h6ac9, 16'h41c4, 16'h2942, 16'h880, 16'h040, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h840, 16'h3164, 16'h5a89, 16'h5a48, 16'h5248, 16'h2123, 16'h820, 16'h213, 16'h840, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h040, 16'h880, 16'h18c1, 16'h2942, 16'h41a4, 16'h72e8, 16'h7b8, 16'h7b8, 16'h93aa, 16'h6aa7, 16'h5a46, 16'h5a26, 16'h5a26, 16'h5226, 16'h5227, 16'h5227, 16'h5a46, 16'h5a46, 16'h5a67, 16'h6aa8, 16'h8bab, 16'h7b4a, 16'h49e5, 16'h1081, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h3984, 16'ha46f, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'ha490, 16'ha490, 16'ha470, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9ce, 16'h9ce, 16'h9ce, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94d, 16'h94d, 16'h93ee, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h8bcd, 16'h8bad, 16'h8bcc, 16'h93ac, 16'h8bac, 16'h8bac, 16'h8bac, 16'h8bac, 16'h8bac, 16'h8bac, 16'h8b8c, 16'h8bac, 16'h8bac, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h838c, 16'h838c, 16'h838c, 16'h838c, 16'h838c, 16'h838c, 16'h838c, 16'h838c, 16'h8b8b, 16'h838b, 16'h836b, 16'h836b, 16'h836b, 16'h836b, 16'h836b, 16'h836b, 16'h732a, 16'h41c5, 16'h20e1, 16'h20e1, 16'h18c1, 16'h18c1, 16'h10a0, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h6288, 16'h62a8, 16'h62a8, 16'h62a8, 16'h62a9, 16'h62a9, 16'h62a8, 16'h62c8, 16'h62c8, 16'h62c9, 16'h6ac9, 16'h6ac9, 16'h6ae8, 16'h6ae9, 16'h6ae9, 16'h6ae9, 16'h73a, 16'h739, 16'h73a, 16'h732a, 16'h7b2a, 16'h7b2a, 16'h7b2a, 16'h72e9, 16'h5a47, 16'h3164, 16'h20e1, 16'h18e1, 16'h880, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h840, 16'h3164, 16'h5a68, 16'h5a48, 16'h5248, 16'h213, 16'h841, 16'h213, 16'h820, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h840, 16'h39a4, 16'h836a, 16'h93cb, 16'h8baa, 16'h8349, 16'h7b49, 16'h8349, 16'h9cb, 16'h6aa7, 16'h5a26, 16'h5a26, 16'h5226, 16'h5226, 16'h5226, 16'h5227, 16'h5226, 16'h5a46, 16'h6266, 16'h6aa8, 16'h8bab, 16'h7b4a, 16'h49c4, 16'h1081, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h840, 16'h3984, 16'ha46f, 16'hacb1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'ha490, 16'ha48f, 16'ha470, 16'ha470, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9ce, 16'h9ce, 16'h94e, 16'h9ce, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94d, 16'h93ed, 16'h93ee, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h8bcd, 16'h8bcc, 16'h8bac, 16'h8bac, 16'h8bac, 16'h8bac, 16'h8bac, 16'h8bac, 16'h8bad, 16'h8bad, 16'h8bac, 16'h8b8c, 16'h8bac, 16'h8bac, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h838c, 16'h838c, 16'h838c, 16'h838c, 16'h838c, 16'h838c, 16'h838b, 16'h838b, 16'h838c, 16'h836c, 16'h836b, 16'h836b, 16'h836b, 16'h836b, 16'h836b, 16'h732a, 16'h41c5, 16'h20e1, 16'h20c1, 16'h20c1, 16'h18c1, 16'h10a1, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h5a88, 16'h62a8, 16'h62a7, 16'h62a8, 16'h62a8, 16'h62a8, 16'h6288, 16'h62a8, 16'h62c8, 16'h62a9, 16'h6ac9, 16'h6ac9, 16'h6ac8, 16'h6ae8, 16'h6ae9, 16'h6ae9, 16'h6ae9, 16'h6ae9, 16'h72e9, 16'h73a, 16'h739, 16'h6ac8, 16'h5227, 16'h41a5, 16'h41c5, 16'h3164, 16'h20e1, 16'h18a1, 16'h860, 16'h020, 16'h020, 16'h020, 16'h020, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h040, 16'h3164, 16'h5a89, 16'h5a48, 16'h5247, 16'h20e3, 16'h861, 16'h2924, 16'h820, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h020, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h00, 16'h00, 16'h020, 16'h5226, 16'h9c2d, 16'h9c2d, 16'h93aa, 16'h8349, 16'h8349, 16'h7b9, 16'ha42c, 16'h6aa7, 16'h5a26, 16'h5a26, 16'h5226, 16'h5226, 16'h5a26, 16'h5226, 16'h5226, 16'h5a46, 16'h6266, 16'h6aa8, 16'h8bab, 16'h7b4a, 16'h41c5, 16'h1081, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h820, 16'h1061, 16'h41a5, 16'ha46f, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hacb0, 16'hac90, 16'ha490, 16'ha490, 16'ha48f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9ce, 16'h9ce, 16'h94e, 16'h9ce, 16'h94e, 16'h94e, 16'h93ee, 16'h94e, 16'h93ee, 16'h93ee, 16'h93ee, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h8bcd, 16'h8bcd, 16'h8bad, 16'h8bad, 16'h8bac, 16'h8bac, 16'h8bac, 16'h8bac, 16'h8bad, 16'h8bac, 16'h8b8c, 16'h8bac, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h838c, 16'h838c, 16'h838c, 16'h838c, 16'h838c, 16'h836c, 16'h836b, 16'h836b, 16'h836c, 16'h836c, 16'h836b, 16'h836b, 16'h836b, 16'h836b, 16'h836b, 16'h732a, 16'h41c5, 16'h20e1, 16'h18c1, 16'h18c1, 16'h18c1, 16'h10a0, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h5a87, 16'h6287, 16'h6288, 16'h62a7, 16'h6288, 16'h62a8, 16'h6288, 16'h62a8, 16'h62a8, 16'h62a8, 16'h62a8, 16'h62c8, 16'h62c8, 16'h62c8, 16'h6ac9, 16'h6ac8, 16'h6aa9, 16'h62a8, 16'h5a67, 16'h5227, 16'h41c5, 16'h3963, 16'h39a4, 16'h41c5, 16'h39c5, 16'h2943, 16'h20e1, 16'h10a1, 16'h840, 16'h020, 16'h020, 16'h00, 16'h020, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h040, 16'h2944, 16'h6289, 16'h5a88, 16'h5247, 16'h18a2, 16'h10a2, 16'h2123, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h040, 16'h840, 16'h861, 16'h10a1, 16'h881, 16'h020, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h820, 16'h526, 16'h9c2d, 16'h9c2c, 16'h93aa, 16'h8349, 16'h8349, 16'h72c8, 16'h9bea, 16'h72a7, 16'h5a26, 16'h5a26, 16'h5a26, 16'h5a26, 16'h5a26, 16'h5226, 16'h5a26, 16'h5a46, 16'h6247, 16'h6a88, 16'h8bab, 16'h7b4a, 16'h49e4, 16'h1081, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h1061, 16'h62a8, 16'h8bac, 16'ha48f, 16'hacd0, 16'hacd0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'hac90, 16'ha490, 16'ha470, 16'ha46f, 16'ha46f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha42f, 16'ha42e, 16'h9c2e, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9ce, 16'h9ce, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94d, 16'h93ee, 16'h93ee, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cc, 16'h8bcd, 16'h93cd, 16'h93cc, 16'h8bcd, 16'h8bcd, 16'h8bad, 16'h8bad, 16'h8bac, 16'h8bac, 16'h8bac, 16'h8bac, 16'h8bac, 16'h8bac, 16'h8bac, 16'h8bac, 16'h8bac, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h838c, 16'h8b8c, 16'h8b8c, 16'h838b, 16'h838c, 16'h838c, 16'h838c, 16'h838c, 16'h836b, 16'h836b, 16'h836c, 16'h836b, 16'h836b, 16'h836b, 16'h836b, 16'h836b, 16'h834b, 16'h73a, 16'h41c5, 16'h20e1, 16'h18c1, 16'h18c1, 16'h18c1, 16'h10a0, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h5a68, 16'h5a68, 16'h6288, 16'h5a87, 16'h6287, 16'h5a88, 16'h6288, 16'h62a8, 16'h62a8, 16'h62a8, 16'h62a8, 16'h62a8, 16'h5aa8, 16'h5267, 16'h4a6, 16'h39a4, 16'h3164, 16'h212, 16'h20e2, 16'h212, 16'h2942, 16'h39a4, 16'h39a4, 16'h3143, 16'h2923, 16'h2943, 16'h211, 16'h10a0, 16'h840, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h040, 16'h2943, 16'h62a9, 16'h6289, 16'h4a27, 16'h1061, 16'h214, 16'h20e3, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h840, 16'h861, 16'h10a1, 16'h212, 16'h2943, 16'h39a4, 16'h39c4, 16'h212, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h49e6, 16'h9c2d, 16'h9c2c, 16'h8baa, 16'h8329, 16'h7b8, 16'h7b8, 16'h93a9, 16'h72a6, 16'h5a26, 16'h5226, 16'h5226, 16'h5a26, 16'h5a26, 16'h5a26, 16'h5a26, 16'h5a26, 16'h6246, 16'h6aa7, 16'h8bab, 16'h7b4a, 16'h49c4, 16'h1881, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h1041, 16'h7b4c, 16'hcdd6, 16'hc573, 16'hb4f1, 16'hacd1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'hac90, 16'ha490, 16'ha48f, 16'ha46f, 16'ha46f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9ce, 16'h9c2e, 16'h9ce, 16'h9ce, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h93ee, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cc, 16'h93cc, 16'h8bcd, 16'h8bad, 16'h8bad, 16'h8bad, 16'h8bac, 16'h8bac, 16'h8bac, 16'h8bac, 16'h8bad, 16'h8bac, 16'h8bac, 16'h8bac, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h8b8c, 16'h838c, 16'h838c, 16'h838c, 16'h838c, 16'h838c, 16'h836b, 16'h836b, 16'h836b, 16'h836b, 16'h836c, 16'h836b, 16'h836b, 16'h836b, 16'h834b, 16'h73a, 16'h41c4, 16'h20e1, 16'h18c1, 16'h18c0, 16'h18c0, 16'h10a0, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h5267, 16'h5a67, 16'h5a67, 16'h5a67, 16'h5a87, 16'h5a88, 16'h5267, 16'h5246, 16'h4a6, 16'h41c5, 16'h39a5, 16'h3184, 16'h2943, 16'h212, 16'h212, 16'h212, 16'h3163, 16'h2922, 16'h2922, 16'h2922, 16'h212, 16'h20e1, 16'h20e2, 16'h292, 16'h2922, 16'h2923, 16'h2922, 16'h18a0, 16'h840, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h020, 16'h2923, 16'h62a9, 16'h5a89, 16'h3185, 16'h861, 16'h3164, 16'h1081, 16'h020, 16'h020, 16'h020, 16'h020, 16'h040, 16'h040, 16'h040, 16'h1081, 16'h213, 16'h2964, 16'h31a5, 16'h39e5, 16'h426, 16'h426, 16'h4a26, 16'h4a6, 16'h212, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h4a6, 16'h9cd, 16'h9cc, 16'h8b8a, 16'h7b28, 16'h72e8, 16'h7b29, 16'h93c9, 16'h72a7, 16'h5a26, 16'h5a26, 16'h5226, 16'h5226, 16'h5226, 16'h5226, 16'h5a26, 16'h5a26, 16'h5a46, 16'h6aa7, 16'h8b8b, 16'h7b4a, 16'h41c5, 16'h18a1, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h020, 16'h020, 16'h020, 16'h020, 16'h840, 16'h62aa, 16'hd617, 16'hde37, 16'hcdd5, 16'hbd33, 16'hb4d1, 16'hacb0, 16'hacb0, 16'hacb0, 16'hac90, 16'hac90, 16'hac90, 16'ha48f, 16'ha48f, 16'ha46f, 16'ha46f, 16'ha46f, 16'ha44f, 16'ha44f, 16'ha44f, 16'ha44e, 16'ha44e, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9ce, 16'h9ce, 16'h9ce, 16'h9ce, 16'h94e, 16'h94e, 16'h94d, 16'h94e, 16'h94e, 16'h94e, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93ed, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h93cd, 16'h8bcd, 16'h8bad, 16'h8bad, 16'h8bad, 16'h8bac, 16'h8bac, 16'h8bac, 16'h8bac, 16'h8bac, 16'h8bac, 16'h8b8c, 16'h8bac, 16'h8b8c, 16'h8b8c, 16'h8b8b, 16'h8b8c, 16'h8b8c, 16'h838c, 16'h838c, 16'h8b8c, 16'h8b6c, 16'h836c, 16'h838c, 16'h838c, 16'h836c, 16'h838b, 16'h836b, 16'h836b, 16'h836b, 16'h836c, 16'h836c, 16'h836b, 16'h836b, 16'h836b, 16'h834b, 16'h73a, 16'h41c4, 16'h20e1, 16'h18c1, 16'h18c0, 16'h18c0, 16'h10a0, 16'h020, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h00, 16'h2945, 
		16'h6b2a, 16'h6b2a, 16'h6ba, 16'h6ba, 16'h62c9, 16'h5a89, 16'h4a27, 16'h3a6, 16'h31c5, 16'h39c5, 16'h39e6, 16'h4227, 16'h4a47, 16'h4a27, 16'h4a26, 16'h39c5, 16'h31a5, 16'h2985, 16'h2985, 16'h2985, 16'h3185, 16'h39a5, 16'h41e6, 16'h4a6, 16'h427, 16'h4a27, 16'h4a26, 16'h39c5, 16'h2964, 16'h2944, 16'h2925, 16'h2925, 16'h2925, 16'h2925, 16'h2945, 16'h2945, 16'h2945, 16'h2945, 16'h2945, 16'h427, 16'h734c, 16'h6bb, 16'h39e7, 16'h427, 16'h4a69, 16'h2945, 16'h2945, 16'h2965, 16'h2964, 16'h2964, 16'h2944, 16'h2944, 16'h2944, 16'h427, 16'h5ac9, 16'h5aca, 16'h62ca, 16'h62ca, 16'h62ca, 16'h62ca, 16'h62ea, 16'h62c9, 16'h427, 16'h2944, 16'h2124, 16'h2124, 16'h2124, 16'h2124, 16'h2124, 16'h2124, 16'h2124, 16'h2945, 16'h62c9, 16'ha48f, 16'ha48f, 16'h9c2d, 16'h93cb, 16'h7b4a, 16'h83ab, 16'ha42c, 16'h836a, 16'h6aea, 16'h6ae9, 16'h6ae9, 16'h6aea, 16'h6aea, 16'h6ae9, 16'h6aea, 16'h6ba, 16'h73a, 16'h7b4b, 16'h9c2e, 16'h8bed, 16'h5aa8, 16'h39a5, 16'h2124, 16'h2124, 16'h2124, 16'h2124, 16'h2124, 16'h2124, 16'h2124, 16'h2925, 16'h2925, 16'h2925, 16'h2925, 16'h2925, 16'h2125, 16'h2945, 16'h2944, 16'h2944, 16'h2945, 16'h6bb, 16'hd617, 16'hde79, 16'hde78, 16'hd637, 16'hc5b5, 16'hbd53, 16'hb532, 16'hb512, 16'hb512, 16'hb512, 16'hb512, 16'hb4f2, 16'hb4f1, 16'hb4f1, 16'hb4f1, 16'hacd1, 16'hb4d1, 16'hb4d1, 16'hacd1, 16'hacd1, 16'hacd1, 16'hacb2, 16'hacb1, 16'hacb1, 16'hacb1, 16'hacb1, 16'ha4b1, 16'ha4b1, 16'ha4b0, 16'ha4b1, 16'ha4b0, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha490, 16'ha470, 16'ha470, 16'ha470, 16'ha46f, 16'h9c70, 16'ha46f, 16'ha46f, 16'ha46f, 16'h9c6f, 16'h9c70, 16'h9c6f, 16'h9c50, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c4f, 16'h9c4f, 16'h9c4f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2f, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h9c2e, 16'h942e, 16'h942f, 16'h9cf, 16'h94f, 16'h94e, 16'h942e, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h94e, 16'h93ee, 16'h8bcd, 16'h5aa8, 16'h39e5, 16'h39e5, 16'h39e5, 16'h39c5, 16'h31a5, 16'h2944, 16'h2124, 16'h2124, 16'h2124, 16'h2124, 16'h2124, 16'h2124, 16'h2124, 16'h2124, 16'h2124, 16'h2124, 16'h2124, 16'h2124, 16'h2124, 16'h2124, 16'h2124, 16'h2124, 16'h2124, 16'h2124, 16'h2124, 16'h2124, 16'h2124, 16'h2124, 16'h2124, 16'h2124, 16'h2124, 16'h2124, 16'h2124, 16'h2124, 16'h2124, 16'h4a69, 
		16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff, 16'hffff
};

	assign width  = 240;
	assign height = 320;

	//assign width  = 239;	for 0 indexed width
	//assign height = 319;	for 0 indexed Height

	assign color  = image[pixel];

endmodule
