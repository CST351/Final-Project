module image(
	input wire [9:0]count,
	output reg [15:0]color
);

reg [15:0] pic[927:0] = '{16'h0000,
16'h001D,
16'h0000,
16'h0020,
16'h0000,
16'h0001,
16'h0010,
16'h0003,
16'h0000,
16'h0080,
16'h0700,
16'h0012,
16'h0B00,
16'h0012,
16'h0B00,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'hF800,
16'h00E0,
16'h0700,
16'h001F,
16'h0000,
16'h0000,
16'h0000,
16'h0042,
16'h4752,
16'h7300,
0000,
0000,
0000,
0000,
0000,
0000,
0000,
0000,
0000,
0000,
0000,
0000,
0000,
0000,
0000,
0000,
0000,
0000,
0000,
0000,
0000,
0000,
0000,
0002,
0000,
0000,
0000,
0000,
0000,
0000,
0000,
00FF,
FFFF,
FFFF,
FFFF,
FFFF,
FFFF,
FFFF,
FFFF,
FFFF,
FFFF,
FFFF,
FFFF,
FFFF,
FFFF,
FF82,
2005,
8247,
D309,
FC47,
D382,
20FF,
FFFF,
FFFF,
FFFF,
FFFF,
FFFF,
FFFF,
FFFF,
FFFF,
FF00,
00FF,
FFFF,
FFFF,
FFFF,
FFFF,
FFFF,
FFFF,
FFFF,
FFFF,
FFFF,
FFFF,
FF82,
2082,
2082,
2082,
2086,
AA09,
FC09,
FC09,
FC82,
20FF,
FFFF,
FFFF,
FFFF,
FFFF,
FFFF,
FFFF,
FFFF,
FFFF,
FF00,
00FF,
FFFF,
FFFF,
FFFF,
FFFF,
FFFF,
FFFF,
FFFF,
FFFF,
FFFF,
FF82,
2047,
D347,
D305,
8282,
2002,
9802,
9802,
9802,
9882,
20FF,
FFFF,
FFFF,
FFFF,
FFFF,
FFFF,
FFFF,
FFFF,
FFFF,
FF00,
00FF,
FFFF,
FFFF,
FFFF,
FFFF,
FFFF,
FFFF,
FFFF,
FFFF,
FFFF,
FF82,
2000,
7000,
7000,
7082,
2009,
FC09,
FC09,
FC09,
FC82,
2082,
20FF,
FFFF,
FFFF,
FFFF,
FFFF,
FFFF,
FFFF,
FFFF,
FF00,
00FF,
FFFF,
FFFF,
FFFF,
FFFF,
FFFF,
FFFF,
FFFF,
FFFF,
FF82,
2082,
2047,
D347,
D382,
209E,
F782,
208F,
738F,
738F,
7382,
2015,
9D82,
20FF,
FFFF,
FFFF,
FFFF,
FFFF,
FFFF,
FFFF,
FF00,
00FF,
FFFF,
FFFF,
FFFF,
FF82,
2082,
2082,
2082,
2082,
2059,
C682,
208F,
7382,
209E,
F746,
D99E,
F782,
2059,
C68F,
7382,
2059,
C682,
20FF,
FFFF,
FFFF,
FFFF,
FFFF,
FFFF,
FFFF,
FF00,
00FF,
FFFF,
FFFF,
FF82,
2086,
D39E,
F79E,
F705,
7282,
2059,
C682,
208F,
7382,
2059,
C646,
D959,
C682,
2059,
C682,
2059,
C646,
D982,
20FF,
FFFF,
FFFF,
FFFF,
FFFF,
FFFF,
FFFF,
FF00,
00FF,
FFFF,
FF82,
2086,
D39E,
F792,
F69E,
F7C5,
A292,
F682,
2059,
C682,
2082,
2046,
D946,
D946,
D982,
208F,
7382,
2059,
C602,
9882,
2082,
2082,
2082,
20FF,
FFFF,
FFFF,
FFFF,
FF00,
00FF,
FFFF,
FF82,
200C,
E592,
F692,
F692,
F692,
F60C,
E582,
2082,
20C6,
B38B,
DC02,
8B9E,
F79E,
F702,
8B8B,
DCC6,
B382,
2082,
20C5,
A205,
7286,
D3C5,
A282,
20FF,
FFFF,
FFFF,
FF00,
00FF,
FFFF,
FF82,
2086,
D392,
F692,
F692,
F692,
F602,
9800,
7082,
2000,
7000,
7000,
7000,
7000,
7000,
7000,
7000,
7082,
2000,
7004,
B886,
D386,
D386,
D382,
20FF,
FFFF,
FFFF,
FF00,
00FF,
FFFF,
FFFF,
FF82,
2046,
D989,
FA46,
D904,
B882,
2082,
2082,
2002,
9889,
FA89,
FA02,
9802,
9889,
FA89,
FA02,
9882,
2082,
2082,
2004,
B886,
D3C5,
A282,
20FF,
FFFF,
FFFF,
FF00,
00FF,
FFFF,
FFFF,
FF82,
20C5,
A286,
D382,
2082,
2015,
9D15,
9D82,
2046,
D902,
9802,
9802,
9802,
9802,
9802,
9846,
D982,
2015,
9D59,
C682,
2082,
2005,
7282,
20FF,
FFFF,
FFFF,
FF00,
00FF,
FFFF,
FFFF,
FFFF,
FF82,
2082,
2059,
C69E,
F746,
D904,
B882,
2002,
9859,
C69E,
F79E,
F79E,
F79E,
F759,
C602,
9882,
2000,
7002,
9859,
C615,
9D82,
20FF,
FFFF,
FFFF,
FFFF,
FF00,
00FF,
FFFF,
FF82,
2082,
2015,
9D9E,
F79E,
F746,
D946,
D902,
9882,
2059,
C682,
2082,
2082,
2082,
2082,
2082,
2059,
C682,
2000,
7004,
B846,
D959,
C659,
C682,
20FF,
FFFF,
FFFF,
FF00,
00FF,
FF82,
2059,
C69E,
F79E,
F789,
FA9E,
F746,
D902,
9882,
2082,
2005,
7286,
D30C,
E592,
F692,
F60C,
E586,
D305,
7282,
2082,
2002,
9804,
B859,
C604,
B815,
9D82,
20FF,
FFFF,
FF00,
00FF,
FFFF,
FF82,
2004,
B846,
D989,
FA46,
D902,
9882,
2005,
72C5,
A286,
D30C,
E592,
F692,
F692,
F692,
F60C,
E586,
D3C5,
A205,
7282,
2000,
7002,
9802,
9800,
7082,
20FF,
FFFF,
FF00,
00FF,
FFFF,
FFFF,
FF82,
2082,
2082,
2082,
2082,
2005,
72C5,
A259,
C605,
72C5,
A292,
F692,
F692,
F692,
F6C5,
A205,
7259,
C6C5,
A205,
7282,
2082,
2082,
2082,
20FF,
FFFF,
FFFF,
FF00,
00FF,
FFFF,
FFFF,
FFFF,
FF82,
2083,
7282,
2082,
20C5,
A2C5,
A29E,
F782,
2005,
720C,
E592,
F692,
F60C,
E582,
2082,
209E,
F7C5,
A2C5,
A282,
2083,
7282,
20FF,
FFFF,
FFFF,
FFFF,
FF00,
00FF,
FFFF,
FFFF,
FFFF,
FF82,
20C6,
B304,
5A82,
20C5,
A205,
729E,
F782,
2082,
200C,
E592,
F692,
F60C,
E582,
2082,
209E,
F705,
72C5,
A282,
20C6,
B3C6,
B382,
20FF,
FFFF,
FFFF,
FF00,
00FF,
FFFF,
FFFF,
FF82,
2083,
728B,
DC83,
7282,
2086,
D382,
2015,
9D82,
2082,
200C,
E592,
F692,
F60C,
E582,
2082,
2015,
9D82,
2082,
2082,
208B,
DC8D,
EDC6,
B382,
20FF,
FFFF,
FF00,
00FF,
FFFF,
FFFF,
FF82,
2002,
8B8D,
ED02,
8B04,
5A86,
D3C5,
A282,
2082,
20C5,
A20C,
E592,
F60C,
E586,
D3C5,
A282,
2082,
2082,
2004,
5A04,
5A83,
728D,
ED8B,
DCC6,
B382,
20FF,
FF00,
00FF,
FFFF,
FFFF,
FF82,
20C6,
B390,
FEC6,
B383,
7204,
5A86,
D30C,
E50C,
E592,
F692,
F60C,
E586,
D304,
5A04,
5A02,
8BC6,
B38B,
DC8B,
DC83,
728B,
DC8B,
DC83,
7282,
2082,
2082,
2000,
00FF,
FFFF,
FFFF,
FF82,
208B,
DC90,
FE8D,
EDC6,
B383,
7204,
5AC5,
A204,
5A86,
D3C5,
A204,
5A04,
5A8B,
DC8B,
DCC6,
B38D,
ED8D,
ED83,
7202,
8B04,
5A04,
5A82,
20FF,
FFFF,
FFFF,
FF00,
00FF,
FF82,
2082,
2082,
20C6,
B390,
FE90,
FE8D,
ED8B,
DC8B,
DC04,
5A8B,
DC04,
5A83,
728B,
DC90,
FE90,
FEC6,
B390,
FE8D,
ED02,
8BC6,
B3C6,
B3C6,
B302,
8B82,
20FF,
FFFF,
FFFF,
FF00,
0082,
2002,
8BC6,
B302,
8B04,
5A8B,
DC90,
FE90,
FE8D,
ED83,
728B,
DCC6,
B302,
8B8D,
ED90,
FE90,
FE8B,
DC90,
FE90,
FE02,
8BC6,
B38B,
DC8B,
DC8B,
DC8B,
DCC6,
B382,
20FF,
FFFF,
FF00,
00FF,
FF82,
2002,
8BC6,
B302,
8B04,
5AC6,
B38B,
DCC6,
B302,
8B8D,
EDC6,
B38D,
ED90,
FE90,
FE8D,
ED90,
FE90,
FEC6,
B38B,
DC8D,
ED90,
FE90,
FE90,
FE8D,
ED8B,
DCC6,
B382,
20FF,
FF00,
00FF,
FFFF,
FF82,
2082,
2004,
5A02,
8B04,
5A04,
5A04,
5A02,
8B8B,
DC8D,
ED90,
FE90,
FE90,
FE90,
FE8B,
DCC6,
B38B,
DC90,
FE90,
FE90,
FE8D,
ED8B,
DCC6,
B382,
2082,
2082,
2082,
2000,
00FF,
FFFF,
FFFF,
FFFF,
FF82,
20C6,
B38D,
ED04,
5A8B,
DC90,
FE02,
8B8B,
DC8D,
ED8D,
ED8B,
DCC6,
B3C6,
B38B,
DC90,
FE90,
FE8D,
ED8B,
DC02,
8B82,
2082,
20FF,
FFFF,
FFFF,
FFFF,
FF00,
00FF,
FFFF,
FFFF,
FFFF,
FF82,
208D,
EDC6,
B304,
5A90,
FE8B,
DC8B,
DC04,
5A83,
7202,
8BC6,
B38B,
DC90,
FE90,
FE8D,
ED8B,
DC02,
8B82,
2082,
20FF,
FFFF,
FFFF,
FFFF,
FFFF,
FFFF,
FF00,
00FF,
FFFF,
FFFF,
FFFF,
FF82,
208B,
DC02,
8B82,
208D,
ED8B,
DC04,
5A82,
20C6,
B38D,
ED8D,
ED8D,
ED8B,
DCC6,
B302,
8B04,
5A82,
20FF,
FFFF,
FFFF,
FFFF,
FFFF,
FFFF,
FFFF,
FFFF,
FF00,
00FF,
FFFF,
FFFF,
FFFF,
FFFF,
FF82,
2082,
20FF,
FF82,
208D,
ED82,
20FF,
FF82,
2002,
8BC6,
B38B,
DC8D,
ED8D,
ED8B,
DCC6,
B302,
8B82,
20FF,
FFFF,
FFFF,
FFFF,
FFFF,
FFFF,
FFFF,
FF00,
00FF,
FFFF,
FFFF,
FFFF,
FFFF,
FF82,
20FF,
FFFF,
FFFF,
FF82,
2082,
20FF,
FFFF,
FF82,
2082,
2082,
2082,
2082,
2082,
2082,
2082,
20FF,
FFFF,
FFFF,
FFFF,
16'hFFFF,
16'hFFFF,
16'hFFFF,
16'hFFFF,
16'hFFFF};

always@(*)
	color = pic[count];
	
	endmodule

	
	
