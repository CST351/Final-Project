//---Example Use---
// GrassTile image1 (
//	.pixel(),
//	.color()
//);

module GrassTile (
	input wire [16:0] pixel,
	output reg [15:0] color
);

	reg [15:0] image [255:0] = '{
		16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h8673, 16'h96b5, 16'h96b5, 16'h8673, 16'h8673, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 
		16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h8673, 16'h8673, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h8673, 16'h96b5, 
		16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h8673, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 
		16'h96b5, 16'haef5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'haef5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'haef5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 
		16'h96b5, 16'haef5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'haef5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 
		16'h96b5, 16'haef5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h8673, 16'h8673, 16'h96b5, 16'h96b5, 
		16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h8673, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h8673, 16'h96b5, 16'h96b5, 
		16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h8673, 16'h8673, 16'h96b5, 
		16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'haef5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h8673, 16'h96b5, 
		16'h8673, 16'h8673, 16'h96b5, 16'h96b5, 16'haef5, 16'h96b5, 16'h8673, 16'h8673, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 
		16'h96b5, 16'h8673, 16'h8673, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h8673, 16'h8673, 16'h96b5, 16'h96b5, 16'h8673, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 
		16'h96b5, 16'h96b5, 16'h8673, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h8673, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'haef5, 16'haef5, 16'h96b5, 
		16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'haef5, 16'haef5, 16'h96b5, 
		16'h96b5, 16'h96b5, 16'h96b5, 16'haef5, 16'haef5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 
		16'h96b5, 16'h96b5, 16'h96b5, 16'haef5, 16'haef5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h8673, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 
		16'h96b5, 16'h8673, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'h96b5, 16'haef5
};

	assign color = image[pixel];

endmodule
